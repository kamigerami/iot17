Kyrkan står mitt i byn .
Det underliga ljudet fick henne upp ur sin säng .
Hon kunde inte komma för hon var sjuk .
Det här vattnet smakar bra .
Jag tycker inte om huset .
Hon är vår granne .
Vi trodde att det var ett flygande tefat .
Detta är huset jag bodde i när jag var barn .
Vi hade roligt på stranden igår .
Jag spelade tennis hela dagen .
De skymtade mannen genom folkmassan .
Han vänjde sig kvickt vid det kalla vädret .
Jag blev tillslut klar med arbetet .
Hon skulle gärna kommit men hon var på semester .
Jag trodde aldrig att ett såhär fint hotell skulle finnas på en sådan här plats .
Detta är deras hus .
Men hon tyckte om barn och gillade sitt jobb .
Hon tycker mycket om att skriva dikter .
Jag kan inte stå ut med detta ljudet längre .
Hon bad mig att se efter hennes bebis medans hon var borta .
Han gnäller alltid på dålig medicinsk behandling .
Stick härifrån , ungjävlar !
Hon är en tillförlitlig person .
Solen skiner .
Den här boken verkar intressant .
Den här boken tillhör skolbiblioteket .
Den här boken handlar om Kina .
Du bör inte lämna barnet ensam .
Studenterna lyssnar på en föreläsning i historia .
Idag mår jag mycket bättre .
Skolan ser ut som en fängelse .
Alla dessa böcker är mina .
Behöver du den här boken ?
Hon ville resa .
Framför oss stod en skrattande flicka .
Han arbetar åtta timmar om dagen .
Jag förstår inte tyska .
Nederländskan är nära besläktad med tyskan .
Många utlänningar pratar bra japanska .
Det är kallt .
Det regnar .
Det är inte viktigt .
Jag minns den första gången .
Det är hett idag .
Kommer du ihåg mig ?
Nu är jag på flygplatsen .
Ingenting saknas .
Föräldrar älskar sina barn .
Jag är väldigt upptagen hemma .
Visa mig ett annat exempel .
Jag har tappat min plånbok .
Igår på morgonen var det väldigt kallt .
Denna stol är ful .
Varför ?
Lycka till .
Vad gör du ?
Vad gjorde du ?
Tack !
Jag ska göra din nya dräkt .
Vilken tid bad han om ditt svar ?
Jag skulle vilja bo i New York .
Han vårdar de gamla fotografierna .
Företaget kämpar för sin överlevnad .
Jag ska fråga honom om det imorgon .
Jag kan inte direkt säga att jag är glad över min pensionering .
Tankfartyget har bara en liten besättning ombord .
Löven ändrar färg i höst .
Skolbarn har förkylningar dubbelt så ofta än vuxna .
Jag orkar inte lyssna mer på hennes klagomål .
Jag ska sluta röka för gott .
Jag erkänner att jag är slarvig .
Jag såg honom igen .
I medicinsk forskning är en av de största problemen att isolera orsaken till sjukdomen .
Han sprang inte tillräckligt fort nog för att hinna med tåget .
Gå in och vinn !
Hur stor summa pengar förbrukar du ?
Det är en vacker Kabuki docka !
Han finslipade en kniv .
Du måste prata med honom angående det
Låt mig fundera ett litet tag .
Hur långt är det härifrån till Hakata ?
Min bror kan springa lika fort som jag kan .
Först och främst måste du leta upp det i ordboken .
Valets resultat kommer snart att bli analyserad .
Han gillar skvaller .
Om ni har något problem så fråga mig om hjälp .
Han blev kry igen .
Han blev en berömd sångare .
I den här tidningen avgränsar jag diskussionen om Emmets ' dyad ' stil i hans verk 1995 .
Han längtar efter att bli en lärare .
Det är underligt för honom att vara borta från skolan .
Han är i en desperat sökning efter fler bevis .
De här blommerna blommar tidigare än vad andra gör .
Den slipsen passar dig tillsammans med din skjorta .
Hon sa att hon inte gillade den , men jag tyckte , personligen , att den var väldigt bra .
Jag ska av nästa station .
Min bil håller på att bli reparerad nu .
Han var sen på grund ut av olyckan .
Ditt motiv var beundransvärt , men inte ditt agerande .
En vis man drar nytta ut av sina mistag .
Han , så som du , är en bra golfspelare .
Förklara hur man tar medicinen är du snäll .
Jag åkte dit med buss och tåg .
Imorgon är det hennes föddelsedag .
Imorgon fyller hon år .
Jag väntade inte länge förän han dök upp .
Kan jag få lite vatten är du snäll ?
Brandmannens ansikte var bistert när han kom ut ur det brinnande huset .
Stilla Havet är det största havet i världen .
Hennes enda önskan var att träffa sin son igen .
Vår lön är liten , fast vi klarar oss .
Jag har varit i mer än tio utländska länder hitills .
Jag sov inte igårnatt .
Jag letar efter ett deltidsjobb .
Du ska få en fin present .
Tack vare Harunas " väder läge " blev Kaoris iver väldigt dämpad .
När måste jag lämna in rapporten ?
Vi måste följa spelets regler .
Ett slagsmål började utan någon anledning mellan dem .
Det är allt jag känner till om honom .
Vet du vad ?
Det är inte den typen av sjukdom som sätter ditt liv i fara .
Han har ett bra rykte som affärsman .
Det är dags att börja röra mig härifrån .
Jag vill att du ska jobba hårdare .
Jösses , vilken oanständig kund !
Eleverna såg alla fram emot sommarlovet .
Han kollade mig rakt i ansiktet .
Jag fick slut på pengar när jag var på besök i Indien .
Jag vet inte vad jag ska säga .
Hon meddelade mig om hennes avfärd .
Det här tyget känns lent .
Han tillgodogjorde det han hade lärt sig .
Det fanns en hatt och en kappa på vägen .
Du kan lika gjärna lämna hemmet på en gång .
Torkan skadade alla skördor där .
Jag kanske gör det ; det beror på omständigheterna för tillfället .
Jag bröt av min tumnagel .
Jag äter upp min hatt om min kandidat inte vinner valet .
Engelska kommer att ta dig en lång tid att bemästra .
På bussar bör ungdomar ge sina sittplatser till de äldre människorna .
Ah , är det så att du blir generad över att bli kallad vid ditt första namn ?
Han flyttade till en varmare plats med omtanke om sin hälsa .
Föraren svängde ratten till höger .
Vad hände ?
Bilen saktar ner .
Nästa koncert kommer att hållas i Juni .
Det hade aldrig slagit henne att han skulle bli bestraffad .
Byron lämnade England för att aldrig komma tillbaks igen .
Min bror måste ha skrivit det här brevet .
Vi talar i Australiens ungdomars vägnar .
Vi är rädda .
Han gifte sig med en vacker flicka .
Varför letar du inte upp det i telefonkatalogen ?
Två andraklassbiljetter till A är du snäll .
Vi vann matchen med 10 mot 4
Jag förklarade det för honom , bara för att förvirra honom .
Det är säkert att han kommer att lyckas .
Vad betyder det ?
Ge mig nyckeln .
Deras trädgård är full ut av väldigt vackra blommor året runt .
Jag hittade en bebis fågel när jag gick i parken .
Han förnekar ingenting för sina barn .
Dom säljer olika saker på den affären .
Han har ett tillräckligt bra omdömde för att inte låna ut pengar till dig .
Läraren var tvungen att utvärdera alla elever .
Segla längst kusten .
Du känner dig ensam , eller hur ?
Låt oss sjunga och dansa .
Den här klänningen skrynklar sig lätt .
Jag vill ha samma ordbok som din syster .
Man ska inte göra sig lustig över andra .
Jag sträckte ut handen mot boken .
Hon ser sin chef som sin far .
John kan inte göra det , och inte jag heller , och inte du heller .
Jag kollade på klockan och visste vilken tid det var .
Vart är den japanska ambassaden ?
Du är bara ung en gång .
Han har redan gått ut .
Jag kommer så fort jag kan .
Man har inte hört något ifrån dom sen dess .
Låna mig din cykel .
Är det öppet på söndag ?
Vi insisiterar på att det skall hållas ett möte så snart som möjligt .
Han var inne i sina egna tanker med handen över hans panna .
Där kommer vår lärare .
Jag tror inte på att det finns någon ond person i denna värld .
Det är skönt och varmt .
Skär köttet i tunna skivor .
Jag vill ha lite pengar .
Han måste köpa en ny cykel åt hans son .
Du har inte den rätta pondusen som chef för avdelningen .
Hur var ditt lov ?
Hur var din semester ?
Vi dekorerade rummet själva .
Jag fick en spark i baken .
Det lilla födelsemärket tog ingenting ifrån hennes skönhet
Vi lagrade höet i stallet .
Det här passet är giltigt för fem år .
Jag har väntat sen klockan sex och det är inte min tur än .
Jag har läst några hundratals böcker .
Om jag visste sanningen skulle jag ha berättat den för dig .
Det var Herr Smith som berättade för mig hur man använde den maskinen .
Jag försökte skriva med min vänstra hand .
En bra lärare måste vara tålmodig med hans elever .
Jag kan inte komma av arbetet nu .
Kan du räkna till tio på kinesiska ?
Koko fortsatte att lära sig fort .
Jag kunde inte förstå något ut av vad han sa .
Rökare sjukskriver sig dubbelt så mycket än vad icke-rökare gör .
Plötsligen förlorade kontorsarbetaren sitt temperament .
Jag visste att han försökte använda pengarna till att bli guvernör .
Vår skola är femton år gammal .
Skicka ditt bagage i förväg .
Jag stod och väntade på en buss .
Vad har du gjort angående reperationen av bilen ?
Oj !
Det är billigt !
Polisen sa till flickorna " Är det här eran bil ? "
När jag väl har blivit vald ska jag göra mitt bästa för er alla som har stöttat mig !
Vi har många jordbävningar i Japan .
Den här datorn är bättre än den .
Tandläkaren drog ut hennes dåliga tand .
Du hade inte behövt köpa ett sådant stort hus .
Jag hoppas att du aldrig blir kommunist .
Vi behöver alla acceptera flödet i dessa tider .
Det ser ut som att det ska börja regna .
Jag är säker på att Teds hostande beror på rökning .
Vi hade det väldigt svårt att hitta busshållplatsen .
Han bor inte där längre .
Jag tappade bort klockan .
Har du varit här sen dess ?
Det här är roten till problemet .
Meg pratar för mycket .
Du kan inte förvänta dig en sådan bra chans igen .
Hennes ansikte blev rött plötsligen .
Tom arbetade hårt bara för att misslyckas på tentan .
Nu finns det ingen återvändo .
Den här firman trycker många läroböcker .
Har far kommit hem ännu ?
Jag tror att jag har råkat på en förkylning .
Han är kortare än Tom .
Vi var fattiga , men glada .
De här reporna syns väldigt mycket så jag skulle vilja få dom reparerade .
Hans uppsats är kopplad till min .
Han köpte den inte i alla fall .
Jag kommer inte att träffa henne igen .
Hon gillar klassiska kompositörer såsom Beethoven och Bach .
Publiken bestod mest ut av elever .
Han har ingen stolthet .
Vi visste inte vilket tåg de skulle vara på .
Vad tycker om Japan ?
Jag önskar dig ett lycka till .
Hela nationen sörjde hjältens död .
Vi är mer eller mindre själviska .
Jag har bott här
Jag fick min son till att träffa doktorn .
Det är dags att du börjar stå på dina två egna fötter .
Jag hoppas att vädret klarnar upp innan vi ger oss av .
Han är oerhört stilig .
Jag kände mig smått illamående .
En kombination av flera misstag ledde till olyckan .
Hon erkände att hon inte kunde prata franska .
Så här långt ser det bra ut .
Det här är året av information , och datorer spelar en ökande viktig roll i vårt vardagliga liv .
Sammanfatta innehållet i 60 engelska ord .
Sluta reta mig .
Ingen dramatiker kan jämföras med Shakespeare .
Hans ilska var förfärlig att se .
Aah !
Min dator frös sig igen .
Kan du förklara hur diskmaskinen fungerar ?
Varför följer du inte med oss till festen ?
Det verkar som att tjuven bröt sig in genom ett fönster på den övre våningen .
Hotellet har en bra utsikt .
Jim kommer inte bra överens med sina klasskamrater .
När jag besökte deras lägenhet var paret precis i ett gräl .
När elden brast ut sov han död som en sten .
Han gjorde äntligen slut med den där kvinnan .
Lite tidigare imorse fick jag ett enanstående nådigt samtal från senator McCain .
Senator McCain kämpade länge och hårt i den här kampanjen .
Och han har kämpat ännu längre och hårdare för det land han älskar .
Han har stått ut med uppoffringar för Amerika som de flesta av oss inte kan föreställa sig .
Det vore bättre om vi var i tjänst framställd ut av denna modiga och osjälviska ledare .
Han svarade inte på mitt brev .
Jag tycker att den sociala sidan är intressant i den nyhetstidningen .
Han är säker på att han kommer vinna matchen .
Vi har ingen snö här .
Hans romaner är för djupa för mig .
Försiktig som han var gjorde han ett oväntat misstag .
Hur många engelska ord kan du ?
Han ägnade all sin tid till att studera historia .
Du kommer inte att finna så många nyheter i dagens nyhetstidning .
Kom hem tidigt , Bill .
De goda nyheterna fick henne att gråta .
Den här pjäsen har ingen humor i sig .
Hästens fall resulterade i ett brutet ben .
Då hade Tyskland en kraftfull armé .
Har du ett recept ?
Vad du har blivit lärd är fel .
Han är lika gammal som jag .
Det fanns inte en själ i sikte .
De är mina bröder .
Far gav mig en veckas veckopeng i förskott .
Far , får får får ?
Nej , får får lamm .
Tomten stod på tomten
Båda föräldrarna lever fortfarande .
De är för nära .
Uppfinnaren är känd över hela världen .
Jag promenerar i skogen varje dag .
Har du någonsin hört talas om Nessie ?
Det var hans anteckningsbok som blev stulen .
Jag måste träffa en tandläkare .
Lägg tillbaks boken där du fann den .
Kärleken kommer så småningomg
Flygfältet på ön är nu täckt med ogräs .
Du måste skörda det du har sått .
Löven virvlade runt i gården .
Jag målade en bild åt dig .
Albert , jag hoppas att du kommer stå vid mig om jag hamnar i problem .
Hon kanske berättade en lögn för mig .
Han gjorde mig en trädocka .
Jag har varit i Paris .
Akiko har några vänner i Frankrike .
Man har funnit olja under Nordsjön .
Han siktade mot fågeln .
Testa den tröjan .
Diska tallrikarna är du snäll .
De har alla självständiga betydelser .
Han klagade över att rätten smakade dåligt .
Vi associerar namnet Einstein med relativitetsteorin .
Jag är nöjd med allt .
Om jag vore en fågel så skulle jag kunna flyga till dig .
Våra eftersträvningar slutade inte med lycka .
Du ska inte tro att det kommer att bli enkelt .
Han vore den sista mannen som skulle göra något sånt .
Han är min chef .
Jag kan inte göra något sånt .
Jag gav det ett försök och tänkte att allting är värt ett försök .
Men att sätta ihop ett sånt här program har jag ingen chans för .
Ett stort djur sprang iväg från zooet .
Skulle du kunna slå in den som en gåva ?
Jag träffade Fred på gatan .
Kom när ni vill .
Regnet föll i mitt ansikte .
De dricker coca-cola .
Mitt uppslagsverk är väldigt användbart .
Armén var tvugna att reterera .
Min mor brukade läsa sagor för mig .
Jag försökte ge henne en gåta .
Även om han säger att han ska återvända till Iran för att gifta sig så är hans planer efter Japan väldigt osäkra .
Han har blivit rundare .
Den gamle mannen och Sjön är en väldigt spännande bok .
Hon fick en stor summa pengar i förskott för hennes nästa roman .
Hon har blivit en helt annan person .
Han var i ett kritiskt tillstånd .
Hon studerade utomlands för att borsta upp hennes engelska .
När lämnar din far hans kontor ?
Jag växlade yen till dollar .
Lärarens elever ser upp till honom .
Du kan alltid räkna med honom i ett nödfall .
Mitt plan går klockan sex .
Läraren kräver utmärkt gjorda arbeten från hans elever .
Skolan ligger en halv mil iväg från mitt hus .
Jag tror att ärligheten kommer att vinna i slutändan .
Han önskar att han kommer besöka Paris .
Rosorna blommar i vår gård .
När kommer du att vara tillbaka ?
Inte underligt att hon inte dök upp för att ge honom ett avsked .
De har gjort slut .
De här verktygen behövs verkligen repareras .
Öppna din mun .
Vem hon är har jag ingen aning om .
En pojke sprang iväg med lite pengar .
Om din chef " plundrar " dig betyder det att du har blivit avskedad .
Kimura joggade i parken varje dag .
Jag undrar om det finns någon mening i att lägga in ordspråk i engelskan ?
Vad är den mest behändliga vägen att ta sig till Tokyo Station ?
Jag höll i festen på egen bekostnad .
Den här gammla bilen går sönder hela tiden .
Det var kallt hela den dagen , och senare började det regna .
Jag är ledsen , vi har inga vaccin .
Ingen kan förneka faktumet att världsekonomin kretsar kring den amerikanska ekonomin .
När brukar du vakna på morgonen ?
Var inte rädd för att göra misstag när ni pratar engelska .
Alla människor andas luft .
Trädgården har blivit proffesionellt anlagd .
I klart väder kan vi se ön härifrån .
Låten var en stor succé .
Det tunga regnet förhindrade mig från att komma ut .
Fotboll är inte nödvändigtvist begränsat till män .
Hon har inte kommit hit än .
Du får inte beté dig så .
Jag åkte ända till London med bil .
Ät mer , annars kommer du inte att få styrka .
Hur länge tar det att gå härifrån till stationen ?
Vi lyckades simma över ån .
En dam , vars man är en känd forskare , kom över från den andra sidan .
Det här huset behöver målas .
Det är dumt av dig att tro på honom .
Det är omöjligt att inte bli fascinerad ut av hans skönhet .
Många barn stannar efter skolan för klubbaktiviteter .
Låt inte din fantasi springa iväg .
Hon kan prata tio språk .
Jag vill veta orsaken till hans frånvaro .
Vi måste kompensera för den förlorade tiden .
Dennis kan göra det fulaste grimasen i staden .
Bortsett från hans häl så var Akilles odödlig .
Antingen har du eller han fel .
Han är före i sin engelska klass .
Matchen blev fördröjd på grund ut av snö .
Han åker skidor i Hokkaido varje vinter .
Arbetet är nu igång .
Hon älskar att se på tennismatcher på TV .
Jag lämnade in ett papper igår .
Hon är en kontorskvinna .
Jag är inte säker på att vi kommer kunna få tag på biljetter ikväll .
Har du någonsin varit i ett främmande land ?
Hans slips matchar bra tillsammans med hans kostym .
Jag kommer inte att glömma bort din vänlighet så länge jag lever .
Det är lite kallt idag .
Vill du följa med ?
Direktörn kontrollerar hans män efter behag .
Isen över ån är för tunn för att kunna bära din vikt .
Solen gör jorden varm och ljus .
Jag hade en väldigt hög feber .
När man är i Rom så gör som romarna gör .
Det här är mina skor och det här är dina .
Färgen av hennes klänning och skor matchade varandra bra .
Han önskade att gud skulle välsigna mig .
Föräldrarna var förtjusta av hennes skönhet .
Lera är en grundläggande ingrediens när man ska göra krukmakeri .
Jag sprang så snabbt jag kunde för att hinna med tåget .
Spiken gick igenom väggen .
Meningar börjar med en stor bokstav .
Det sägs att han är född i Afrika .
Det är söndag imorgon .
Ingen väntar vid busshållplatsen .
Vi kanske har missat bussen .
Grekerna äter också ofta fisk .
Vi misslyckas att förstå ordets mening .
Hon slöt in det i papper .
Ring mig klockan fyra .
Jag måste ta det första tåget .
Han var inte samma glada man han en gång var .
Verkligen .
What kan jag göra ?
Vi såg båten gungande ute på den stormiga sjön .
Jag behöver inte din hjälp .
Hur länge kommer du att vara i Japan ?
De seglade runt världen .
Han är medveten om hans eget fel .
Stunden kommer att komma då du känner dig skyldig för det .
Jag känner mig inte för att träffa henne nu .
Han sprang för fort för att vi skulle kunna hinna ikapp .
Olyckan skedde i det hörnet .
Han är ofta förskenad till skolan .
Du är den sista personen jag förväntade mig att träffa här .
Den här dramaserien kommer att sändas imorgon .
Människorna skrattade tills hon sa " Brinn ! " .
Du är väl inte rädd för spöken ?
Medicinen smakar beskt .
Skulle du vilja följa med på en promenad ?
Hon lever ett olyckligt liv .
Jag är hungrig .
Jag är hungrig för jag har inte ätit lunch .
Jag tror inte att det kommer att regna i morgon .
Jag är bäst .
Ärligt talat , hans tal är alltid tråkiga .
Han stal plånboken av mig .
Mina pengar är slut .
Tack för din förklaring .
Vad ?
Jag pratar inte japanska .
Jag kan inte japanska .
Vad kostar det ?
Jag förstår inte .
Vad är det ?
Vad består aspirin av ?
Sluta fråga mig om en drink !
Gå och hämta en själv .
Vad skulle världen vara utan kvinnor ?
Du kan inte prata så högt här .
Det är för mörkt för att jag ska kunna läsa .
Du får inte parkera bilen på denna gata .
John och Mary har känt varandra sedan 1976 .
Nancy , här är ett brev till dig .
Hon är inte så ung som hon ser ut .
Denna blomma är gul , men alla de andra är blåa .
Jag tror att han var arg .
Mörker är frånvaro av ljus .
Vems cykel är det här ?
Ett , tre och fem är udda tal .
Min fru hatar katter .
Det här gamla bordet används fortfarande .
Han gillar att sjunga populära sånger .
Jag har fullt upp just nu .
Alla hästar är djur , men inte alla djur är hästar .
Jag gillade henne inte till en början , men nu gör jag det .
Du måste vara på stationen senast klockan fem .
Hon är en duktig tennisspelare .
Nederländerna är ett litet land .
Tecknet visar att svaret är rätt .
Läkaren bad herr Smith om att sluta röka .
Bryt chokladen i små bitar .
En gammal man vilade sig i skuggan av trädet .
Jag visste inte när jag skulle slå av maskinen .
Man skall älska sin mor .
Ge mig lite vatten , och det snabbt .
Jag är väldigt glad att se dig igen .
De gav oss jobben .
Vi är bjudna på middag .
Det är ganska kallt .
Det överraskar mig inte .
Det där är inte en kniv .
Det HÄR är en kniv !
Han älskade att resa .
En dag fann jag en bok där .
En gång fann jag en bok där .
Kan du visa mig vad du har köpt ?
Dessa två bröder liknar varandra .
Vi ska mötas på stationen klockan nio .
Var snäll och vänta i fem minuter .
Ta det inte personligt .
Han hade tänkt att gifta sig med henne .
Denna skrivmaskin har använts mycket .
Bilden hänger upp och ned .
Jeg vet inte om han kommer att besöka oss nästa söndag .
Jag är från Tokyo , Japan .
Hur är det ?
Jag har inte sett dig på evigheter !
Det är två elever borta idag .
Jag blir ofta förväxlad med min bror .
Klimatet är behagligt .
Jag började tillsammans med två resande kompanjoner .
Du kan lita på honom .
Han tror fortfarande på hennes ord .
Företaget gick i konkurs .
De är väldigt intresserade av astronomi .
Han är en poet .
Vilket tåg tänker du ta ?
Brevets innehåll var hemligt .
Han är stolt över att ha tagit examen vid Tokyo Universitet .
De har ingen annanstans att gå .
De har ingen annanstans att ta vägen .
Jag älskar dig .
Allt som är för dumt för att sägas sjungs .
Jag hittade en lösning , men jag hittade den så fort att det inte kan vara den rätta .
Han har faktiskt inte ätit kaviar .
Bjud oss på middag på restaurang !
Min pappa promenerar varje dag .
Cuzco är en av de intressantaste platserna i världen .
De som inte önskar gå behöver inte det .
Han visade mig sin frimärkssamling .
Det här stället har en mystisk atmosfär .
Vi såg barnet kliva på bussen .
Jag har en katt och en hund .
Katten är svart och hunden är vit .
Gillar du golf ?
Jag känner tjejen som spelar tennis .
" Jag är hungrig " , sa den lilla vita kaninen , så de stannade och åt blomman av en stor hyasint .
Folk säger ofta att japanska är ett svårt språk .
Folk säger att han aldrig dör .
Vi ses !
Om han hade tagit mina råd så hade han varit rik nu .
Han började lära sig spanska genom radion .
Jag förväntar mig en tunnelbanestation här i framtiden .
Jag har inte hört något från honom sen dess .
Jag känner på mig att han känner till hemligheten .
Jag var född och uppfostrad i Matsuyama .
Lejonet öppnade sin enorma mun och vrålade .
Hon rynkade pannan .
Det är en självklarhet att grundläggande mänskliga rättigheter bör respekteras .
Amen ge dig iväg .
Påminn att posta breven är du snäll .
Hur stor är New York Citys befolkning ?
Glada är de som känner till värdet av hälsa .
Den här målrätten är lämplig för tre .
Vi gör det när han kommer .
De plaskade vatten i mitt ansikte .
Företaget bidrar med sjukvård och livförsäkringar åt alla dess anställda .
Inget är så hemskt som en jordbävning .
Det händer att dörren är öppen ibland .
Det tjänar inget till att bråka med honom om det .
Hans bil kolliderade med ett tåg .
Precis när hon skulle lämna affären så såg hon en vacker klänning i fönstret .
Jag vill köra ett Windows 95 spel .
Jag gillar engelska , men jag är inte så bra på att tala det .
Stormen utbrast .
Nej , hon har aldrig blivit förälskad .
Jag betalar notan .
Kommer hon med ?
Var rädd om dina möten med andra för du vet aldrig om du bara möter personen en gång om livet .
Hon frågade mig om jag mådde bra .
Men jag kan aldrig hålla mig .
Hur långt kommer det att ta för att bli återställd ?
Jag såg henne på festen .
Det kan inte vara sant .
En man kan leva och vara frisk utan att döda djur för mat .
Därför deltar han i att ta djurs liv enbart på grund ut av hans aptit om han äter kött , och att bete sig så är omoraliskt .
Han är ostoppbar just nu men frågan är hur länge han kan hålla sig kvar vid sin höjdpunkt ut av sin karriär .
Den här vägen kommer att leda dig till parken .
Säg vad vi ska göra härnäst .
Molnigt med återkommande regn .
Har du gjort klart din engelska läxa än ?
Med små steg började rosbuskens knoppar blomma .
Det kommer att regna den här eftermiddagen .
Vi lekte ofta mamma pappa barn i parken .
Någon verkar ropa på mig .
En revolution bröt ut i det landet .
Fattig som hon var gav hon honom det lilla hon hade ut av sina pengar .
Domaren utgav honom som vinnare .
Den räven måste ha dödat hönan .
Jag kan inte förstå alls vad det är du säger .
En bebis är inkapabel ut av att ta hand om sig själv .
Han sov gott igårnatt .
Vilken typ av sport gillar du ?
Hon måste ha varit väldigt vacker när hon var ung .
I amerikansk fotboll har försvaret en specifik roll .
När gick du upp imorse ?
Tallriken slank från hennes hand och krashade ner i golvet .
Först och främst måste vi bestämma oss för ett namn .
Jag har inga pengar .
Det är en bild som jag gillar väldigt mycket .
Lucy är en fin liten flicka .
Känner du till någon doktor som kan prata japanska ?
De här skorna är en aning för stora .
De här skorna sitter inte särskilt bra .
Det stämmer att projektet är en svår uppgift , men herr Hara kommer att kunna göra det .
Han bor på andra sidan floden .
Staten New York är nästan lika stort som Grekland .
Lägg till vatten och blanda ihop det till en mjuk deg .
Du har friheten att använda detta rum hur du än vill .
För Amerikaner , på andra sidan , är det mer troligt att ta risker i hopp om att uppnå stora framgångar .
Jag är inte mannen som du en gång kännde mig som .
Han lämnar alltid sina verk gjorda till hälften .
Helen håller alltid sitt rum rent .
Solen går upp i öst och ner i väst .
Han skickade mig ett föddelsedagskort .
Till hennes sorg hade hennes son lämnat henne ensam .
Jag kännde igen henne stunden jag såg henne .
När jag tänker på de där eleverna får jag huvudverk .
Han gick inte , och det gjorde inte jag heller .
Skulle du kunna säga mig vilken station som ligger närmast ditt arbete är du snäll .
Han svarade genom att ge " OK " gesten .
Den nya maskinen kommer att ta upp en massa utrymme .
Vi gick på picnic till kullen .
Inget sött utan svett .
Men snart skulle han inte kunna gå , skriva eller ens äta själv .
Kom snälla du , jag är ivrig över att se dig .
Den här låten påminner mig alltid om mina skoldagar .
En dator är inte mer levande än vad en klocka är .
Min bror vågade ej att simma över floden .
Jag brukade åka skidor på vintrarna .
Pojken som bor här intill kommer ofta hem sent .
Hon brann med svartsjuka .
Har du gjort något nyårslöfte ?
Stålproduktion nådde uppskattat 100 miljoner ton förra året .
Vi får se vad som händer .
Mannen som jag besökte var Mr Doi .
Lyssna noga är du snäll .
Han har gjort sitt yttersta för mig .
Jane ska undervisa våra elever från och med nästa vecka .
Hon är sig själv igen .
Han drog förbi en vän .
Det är en fots längd mellan de två husen .
Missförstå mig ej , vi gör inga löften .
Jag har bestämmt mig för att vara glad för det är bra för min hälsa .
En helicopter åkte runt över oss .
Nöjet av att resa runt är vanligt hos nästan alla personer .
Ann kommer inte till våran fest .
Han blev nästan dränkt .
Jag är inte trött alls .
Att föra en dagbok är en bra vana .
Vi prövar en helt ny metod .
När hennes grannar var sjuka frågade hon doktorerna att ge dem medicinska hjälpmedel .
Min son som går i femteklass har förflyttat sig till skolan i Nagoya från Shizuoka .
Han har gått till Nagoya för affärer .
Tvål har förmågan att få bort smuts .
Virvelvinden tog med sig förlust av regn till det distriktet .
Han sa att han hade köpt den boken där dagen innan .
Jag tenderar till att dra till mig förkylningar .
Det är en bra regel varsomhelst att se åt båda håll innan du gå över gatan .
Det här är den vackraste utsikten som jag någonsin sett .
Hon kan prata både engelska och tyska .
Han stannade hos hans fasters hus
Han stannade hos hans mosters hus .
Han sov över hos hans fasters hus .
Han sov över hos hans mosters hus .
Jag skaffade en ny högtalare i den affären .
Håll käften , eller så slår jag ner dig .
Att träna varje dag är nödvändig för din hälsa .
Jag har en känsla på mig att hon kommer att komma idag .
Du är riktigt klusmig av dig va !
Vårt lov kommer snart att nå sitt slut .
Det är bara ett par få minuter kvar tills tåget går och hon har inte dykt upp än !
Min mormor blev åttioåtta år gammal .
Vad skulle hända om han skulle komma försent ?
Tack vare televisionen är pojkar och flickor benägna att ej läsa böcker .
Kämpa !
En katt dök upp från baksidan av drapperiet .
Kastrullen kokar .
Deras nationalism var en ut av orsakerna till kriget .
Han är ivrig över att tillfredställa allihop .
Tog du ett bad ?
Jag kommer att kunna träffa honom nästa år .
Han fuskade under provet genom att kopiera från flickan framför honom .
Du är lyckligt lottad som har sådana vänner .
Priset på olika maträtter varierar från vecka till vecka .
Vare sig du lyckas eller inte beror på dina egna ansträngningar .
Flickan var alldelles utom av sig av sorg .
Det brukade finnas en restaurang framför den här busstationen .
Hon var nära på att drunkna .
Jag kanske har lagt den på bordet .
Han har bara en tröja för resten av dom är på tvätt .
Klockan är redan elva .
Det är dags att du kommer i sängs .
Den gamle mannen var inte så elak som han såg ut att vara .
Jag tog det förgivet att hon skulle hålla med mig .
Herr Crouch , vad gör du ?
Det var inte förrän igår jag fick nyheterna .
Tåget var fullt med passagerare .
Kan du finna den ?
Kan du hitta den ?
Det tog honom tio minuter att lösa problemet .
Jag läste brevet åt honom .
Han ansträngde sig ej .
Det är nödvändigt för oss att sova gott .
Kvinnan som sitter där borta är hans nuvarande fru .
De passar varandra på grund ut av deras närliggande intressen .
Avdokaten insisterade över klientens oskyldighet .
Jag vill komma ut härifrån !
Han är väldigt upptagen med att skriva till hans vänner .
Det är nödvändigt att bekämpa AIDS med vilket vapen vi nu än behöver !
Det började regna kraftigt för mer än tre timmar sedan .
Han försökte hårt i förgäves .
Vad hände på bussen ?
När kom demokrati in i existens ?
Har du hört honom sjunga ?
Vad menar du med " den " ?
Jag har problem med att pulvermedicin .
För vilken anledning bröt du dig in i huset ?
Hon instämmde med våra begär .
Min rygg gör fortfarande ont .
Möt konsekvenserna .
Åker den här bussen till Park Ridge ?
John ' s mor ser så ung ut så att hon ofta misstas för en ut av hans äldre systrar .
Han är bra på att imitera hennes irländska brytning .
Banken tar hand om pengar åt folk .
Hur stor är han ?
Hur gammal är han ?
Han högg av en gren från trädet .
De stack vid klockan 5 , så de borde vara hemma vid 6 .
Jag råkade höra konversationen .
De skillde sig förra året .
Han förklarade hans situation för mig .
Kommer du att lyckas med att reparera min bil ?
Det är tyst här om nätterna .
Det börjar bli molnigt .
Det kanske börjar regna snart .
Även om jag var trött så försökte jag mitt bästa .
Han var arg över att jag hade kränkt honom .
Det här är ett sådant enkelt problem så att vilken elev som helst kan lösa det .
Provresultatet visade hur mycket han hade pluggat .
Hur sent kan jag ringa ?
Man lär sig ut av erfarenheter .
Vi kan inte leva utan luft .
Jag kanske skriver ett brev åt dig .
Även fast jag satt i solen så kände jag mig kall .
Dina framgångar beror på dina ansträngningar .
Jag tycker inte om att handla varje dag men jag måste göra det .
Det är ingen idé att prata med honom .
Han lyssnar aldrig .
Vad ska du ha ?
Mars är desto mer intressant för dess närliggande likhet med vår jord .
Kom hit om två veckor från och med idag är du snäll .
Jag fruktar det .
Han har tre familjemedlemmar att försörja .
Tom förlöjlar sig alltid över John på grund ut av hans dialekt .
Tom gör alltid narr ut av John på grund ut av hans dialekt .
Han ägnade sig helt helhjärtat åt henne .
De smyckrade upp rummet med blommor .
" Är drinkarna gratis ? "
" Bara åt damer . "
Jag tror att han är en schyst kille .
Tack för att du tog mig hit .
Han kände sig fram genom mörkret .
Vi behöver tänka över problemet mer försiktigt .
Tiden är mogen för en drastisk förändring .
Båda eleverna klarade av alla prov .
Jag minns mannens ansikte men jag kommer ej ihåg hans namn .
Jag representerade mitt universitet på konferansen .
Hon var snäll och tog mig till sjukhuset .
Jag har klättrat upp för berget Aso .
Dina föräldrar kom inte , eller hur ?
Hon lämnade scenen förra året .
Jag vet inte om jag har tid att göra det .
Jag gillar varken den ena eller den andra kakan .
Vi måste dra tillsammans och supa någon gång .
Hon försökte hoppa upp en andra gång .
Jag avbröt min hotelreservation .
Vi har väldigt besvikna över att höra nyheterna .
Förlåt , men jag hör dig ej så bra .
" Om det är pengar så lånar jag inte ut något " sa jag kort och gott .
Finns det något vatten i kannan ?
Om jag blir rik så kommer jag att köpa den .
Nancy handlade lite på vägen .
Hej Mimi !
Hur mår du ?
Gör det som du tycker är rätt .
Han drog sig tillbaks till sitt rum efter kvällsmaten .
Jag sa till henne att kvickt göra klart rapporten .
Va ?
Vad falls ?
Ska de inte använda sig ut av mitt förslag ?
Han är känd som den bäst advokaten i den här staden .
Allt du behöver göra är att berätta sanningen .
Hans affär orsakade stora förluster .
Det är just den boken som jag har väntat så länge på för att läsa .
Skulpturerna är av högt värde .
I Japan behöver vi sätta på ett sextiotvåyenfrimärke på ett brev .
Vi körde för snabbt för att njuta ut av det vacka landskapet .
Jag var missnöjd över att det fanns så lite att göra .
Han hade en underlig dröm .
Jag har redan gjort det .
Han var mer än en kung .
Jag ska ringa om det imorgon .
Jane spelade väl inte tennis ?
Jag såg mig omkring men fann ingenting .
Enligt många religioner är äktenskapsbrott ett brott .
En man vars fru är död kallas för en änkling .
Var inte dum .
Franska talas i en del av Kanada .
Vi tipsade dom om att börja tidigt .
Hans mål är att bli en lärare .
Våg efter våg forsade upp på stranden .
Det tog henne hela eftermiddagen att göra klart arbetet .
Han gör vin av grapefrukt .
Hur långt ifrån ligger nästa bensinstation ?
Direktören gav exakt det svaret som jag letade efter .
Den här rörelsen från landbygds- till stadsområden har pågåtts i över tvåhundra år .
Jag trodde att han var en doktor .
Det är upp till dig .
Han sjöng en sång .
När vi kom hem hade solen gått ner helt och hållet .
Kan du säga till mig när jag ska av ?
Hon skrek i sin förvåning .
Mormor bar bordet själv .
Farmor bar bordet själv .
Är hon gift ?
Hej !
Hur mår du ?
En handfull datorer stals vid inbrottet .
Mig vantar kort .
Alla människor äro födda fria och lika i värde och rättigheter .
De äro utrustade med förnuft och samvete och böra handla gentemot varandra i en anda av broderskap .
Ja .
Sonen ställde en fråga till hans mor .
Var såg du henne ?
Oljuden väckte mig .
Fundera på det .
Jag kan inte Svenska .
Jag ska köpa en bil .
Igår hon köpte grönsaker .
Är han en läkare ?
Jag brukar inte dricka kaffe utan socker .
Jag vet inte .
Vad gör han nu ?
Är du upptagen ?
Akiko har flera vänner i Frankrike .
Vad har du i din påse ?
Tack så mycket !
Jag vet inte precis när jag ska vara tillbaka .
Han bor med sin föräldrar .
Han har skrivit en bok om Kina .
Vi behöver en ambulans .
Hatten är din .
Han borde avslöja alltihop och möta konsekvenserna .
Ingen ut av eleverna var försenade till skolan .
Flickan gick in i rummet .
Kom så skakar vi mattan .
För träd är grenar vad lemmar är för oss .
Hur många minuter blir det om du omvandlar 48 timmar till minuter ?
Jag skulle vilja ha en till kopp kaffe .
Vi ska ha prov i engelska imorgon .
Strax innan bröllopet skrek den berusade fadern : " Jag kommer inte att lämna ut min dotter till någon främling ! " till brudgummen .
Han tycker om att se på TV .
Det här halsbandet som tillhör Jane är en gåva från hennes mormor .
Det här halsbandet som tillhör Jane är en gåva från hennes farmor .
Jag vill inte ha den längre .
Jag skulle vilja äta äpple paj .
Han är i tjänst inatt .
Den här sången är en kärlekssång .
Är det en ko eller bisonoxe ?
Mötet sköts upp tills nästa fredag .
Finns det någon som kan uttala det här ordet ?
Jag började att läsa boken .
Hur anmäler jag en stöld ?
Var snäll mot henne , Bill .
Min fars bil är gjord i Italien .
Om du strular till det så kan det inte göras om , så strula inte till det !
Det enda gången då folk inte tycker om skvaller är när du skvallrar om någonting om dem .
Huset brinner .
Han kan varken läsa eller skriva .
Market Square är det historiska centret i staden .
Senaste gången var det en naturlig födelse .
Utan vatten så skulle vi snart dö .
Är du allergisk mot någon medicin ?
Jag vill att du läser det här engelska brevet .
Jag förstår exakt hur du känner dig .
Ditt hus är tre gånger så stort än mitt .
Det verkade som om hon redan hade fått pengarna .
Senatorn anklagade mig för att ha förvrängt datan .
Jag fick ett brev som informerade mig om hans ankomst .
Vem är det som bor här intill ?
Han är en munter kamrat .
Jag antar att du beredd på att ta risken .
Du ser blek ut .
Du måste gå vare sig du gillar det eller ej .
De gifter sig nästa månad .
" Har inte vi träffas någon gång ? " frågade eleven .
Ingen kan lyckas med något utan ansträngning .
Jag kom enbart för att ge besked om faktumet .
Jag vet inte vad det är .
Han kan inte alls engelska .
Jack kan engelska .
En flicka ringde mig .
Var är Britney Spears ?
Jag skriver til Erwan Le Bourdonnec .
Vilken färg är din hår ?
Han borde inte komma tillbaka här .
Det är flickan som jag känner väl .
Jag kan sjunga det på engelska .
Vi har för många lektioner .
Är det din bok , Mike ?
Jag gillar att läsa deckaren .
Jag vil inte ha en smörgås .
Ska han dö ?
Vi behöver pengar .
Dina skor är här .
Frukost är en smörgåsbord .
Få jag låna din bil ?
Är du inte trött ?
Jag har ingen pengar .
Bob är min vän .
Kom och drick té med mig .
Det tog nätt och jämnt en timme .
Vad skulle du vilja äta ?
Jag har två bröder .
Kan hon franska ?
Hej .
Jag heter Farshad .
Skytten dödade hjorten .
Hon gav honom en klocka .
Jag är arbetslös .
Jag valde fel flagga på grund av ett missförstånd .
Jag älskar dig mer än du älskar mig .
Grattis på födelsedagen !
Dessa tvillingbröder är lika som bär .
Det är mycket ovanligare för en person att vara politiskt medveten än att vara politiskt aktiv .
Det är för att jag ska höra din röst ordentligt .
Jag har lite pengar .
Det regnade igår .
Det förvånar mig inte .
Plastfolie är tillverkad i polyethylen .
Du berättar inte sanningen .
Vad man icke kan tala om , därom måste man tiga .
Jag har en svår smärta i ryggen .
Vet du inte att han gick bort för två år sedan ?
Jag vill ha ett eget rum .
Morötter och rovor är ätbara rötter .
Jag gick hemifrån vid sju .
Du kan lämna rummet nu .
Han gav oss kläder , och pengar också .
Liftarna var närapå förfrusna när de hittades .
Du kan använda ett lexikon till den här tentamen .
Han har en plats i parlamentet .
Hans utställning på stadsmuséet tilltalade mig inte alls .
Om det var han så kunde han gjort sämre ifrån sig .
Jag kommer att åka oavsett väder .
Han kommer inte att misslyckas vid examinationen .
Huset höll på att målas av min far .
Det är bara en dröm .
De vann faktiskt .
Sedan jag återhämtade mig från min allvarliga sjukdom ter sig hela skapelsen vacker för mig .
Kan jag avboka den här biljetten ?
Tårar föll från hennes ögon .
I framtiden vill jag bli en TV-presentatör .
Tanken på att hon skulle möta den berömda sångaren fick henne att rysa av spänning .
Du kan använda mitt skrivbord om du vill .
Han utförde arbetet så gott han förmådde .
Förespråkare av ökade importavgifter är oense med varandra .
Han stannade upp mitt sitt anförande .
Är du för eller mot det här ?
Jane är fet , ohövlig och röker för mycket .
Men Ken tycker att hon är förtjusande och härlig .
Det är därför de säger att kärleken är blind .
Jag är rädd att jag inte kommer att vara ledig förrän examinationen är slut .
Polisen hann ifatt honom .
Jag är ledsen , vi har helt slut på manti .
Städa rummet .
De säger att han har varit död i två år .
Min bror är intresserad av det man kallar popmusik .
Mitt armbandsur behöver lagas .
Jag håller inte med din åsikt .
Jag håller inte med dig .
Din fråga hör inte till ämnet .
Paula måste hjälpa hennes pappa i köket .
Vår telefon fungerar inte längre .
Jag skulle behöva laga den .
Jag tycker att det är ganska konstigt att han inte skulle veta någonting sådant .
Vi ska ha barn .
Jag äter här .
Nu behövs inte bara ord , utan också handling .
Jag har en bok om fiske .
Låt oss göra det någon annan gång .
Det är bara en ursäkt .
Min bror har aldrig bestigit Mt Fuji .
Jag är mycket hungrig .
Jag är jättehungrig .
Du med , min son !
Jag skapade en genväg på skrivbordet .
Jag heter Jack .
Ett ögonblicks tvekan kan kosta en pilot livet .
Jag visste inte hur jag skulle svara på hans fråga .
Jag älskar min mamma .
Han är en gentleman .
Jag är från Kyoto .
Hur skulle det vara med en kopp te ?
Ge mig en kopp te , är ni snäll .
Min mor tycker mycket om té .
Klockan är tio i åtta på morgonen .
Han gav mig kaffe trots att jag hade bett om té .
Lite mer mjölk i kaffet , tack .
Jag föredrar kaffe framför té .
Isen smälter .
Ge mig lite mer té .
Skulle ni vilja ha en kopp té ?
Beatles bestod av fyra musiker .
Vill ni ha té eller kaffe ?
Flickan höll på att koka te till åt sin kamrat .
Jag bad honom att koka lite té .
Han bor i Kyoto .
Hon bor i Kyoto .
Ena sidan av ett mynt kallas för ' krona ' och den andra kallas för ' klave ' .
Fler säljer snus med stavfel .
Om du har ett problem med råttor och möss , så kan du skrämma dem med ultraljud .
En man hotade hiv-smitta två sjuksköterskor .
Jag väcks av ljudet från vågorna .
De känns ovanligt nära , och det är de också .
Tjuven bröt upp fönstret .
Koka lite vatten .
Kan du tillaga det här köttet lite mer ?
Jag orkar inte mer !
Jag har inte sovit på tre dagar !
Det kommer att regna .
Han har kanske många flickvänner .
Hon låtsades att hon inte hade hört vad jag sa .
Vi kan se tusentals stjärnor på himlen .
Jag arbetar 3 timmar varje söndagsmorgon .
Färglösa gröna idéer sover rasande .
Hur gammal är du egentligen ?
Hur gammal är du ?
" Hur gammal är du ? "
" Jag är sexton år . "
John er mun hærri en Mary .
Jag heter Hopkins .
Det är något med honom som jag inte gillar .
Skulle du kunna skriva ner länken till den sajten ?
De gick tidigt .
Jag minns när Anna berättade att hon blivit kär .
Körd rimmar på skörd .
Jag anbefaller dig åt Gud .
Vi bygger landet i gärning och ord .
Om du har följt vad jag skrivit tidigare .
Hur många studerade på medeltidens universitet ?
Han kände sig trött .
Flygplanet ankommer klockan åtta .
Jag har inte berättat för mormor om städhjälpen .
Allan har lämnat oss .
Honom har hon inte sett på länge .
Vi frågade honom vad han hette .
Jag har precis kommit tillbaka från Sverige .
Förstår ni vad hon menade ?
Vi vill inte vänta längre .
Huset ligger vackert till .
Föraren körde om bilen .
Hon blev polis .
Jag tycker inte om honom , men jag gillar henne .
Jag måste gå nu .
Hon hade inte råd .
Han målar inte väggarna utan tapetserar dem .
Skål !
Vill du äta ?
När kommer han ?
Vem är du ?
Har du barn ?
Vill du gå ?
God dag .
Detta är ett litet steg för en människa men ett jättekliv för mänskligheten .
Var arbetar du ?
Det här är en turkisk tradition .
Den här är ny .
Jag vill inte bo ensam .
Ursäkta att du fick vänta länge .
Vet du inte vad som hände igår ?
Jag vet inte när mor kommer hem .
Ta din sudd och sudda bort dessa tecken .
Är du japan ?
Vi gick i samma klass på högstadiet / gymnasiet .
Jag har inte sett honom på några år .
Berätta för mig när du ger dig av .
Jag vill dricka en kopp kaffe .
Detta är fakta .
Hon gillar inte fotboll .
Jag är upptagen , så jag kan inte gå .
Vårt skolbibliotek är väldigt litet , men det är nytt .
Slips passar dig .
Du passar i slips .
Slipsen och min kavaj matchar inte .
Om jag är homosexuell , är det en synd ?
Jag har ett par skor .
Jag kommer genast hem .
Det är hennes födelsedag imorgon .
I morgon är det hennes födelsedag .
Hon är intelligent .
Du är verkligen jättebra .
Godmorgon , Mike .
Öppna flaskan , tack .
Välj en person , tack .
Vi förbereder oss för att gå ut .
Jag känner kvinnorna där .
Dagarna blir längre och längre .
Min pappa har åkt för att fiska .
I så fall tror jag att du bör komma idag .
Gillar du fisk ?
Vad sägs om den här röda mössan ?
Fram tills nu har de jobbat mycket hårt .
Är du nöjd med ditt nya hus ?
Vad gjorde Kumi ?
Min bil är i din tjänst .
Helsingfors är huvudstaden i Finland .
Hon hade hjärtformade örhängen .
Kan du vara snäll och vänta en minut ?
Jag har många vänner som hjälper mig .
Jag måste gå och sova .
Jag har ingen katt .
Det här äpplet är väldigt rött .
Svara på frågan .
Vilken är din gitarr ?
Stillhet är guld .
Varför är du så ledsen ?
Ska du äta hemma eller ute ?
Vem har skrivit denna bok ?
Han är nöjd med sitt jobb .
New York är en stor stad .
Coles axiom : Summan av intelligensen på planeten är en konstant ; befolkningen växer .
Jag är törstig .
Hoppas medan du lever !
Det tog dem två år att bygga huset .
Vilket djur gillar du mest ?
Hans förklaring var inte tillräcklig .
Han övertalade sin fru att inte skilja sig .
Jag älskar att resa .
Vi är säkra på vår vinst .
Jag förlorade medvetandet .
Du borde skriva om denna mening .
Tom hittar alltid fel hos henne .
Har du inte bestämt dig än ?
Han brast ut i gråt .
Den andra fungerar inte .
Du var hemma i går , inte sant ?
I dag mår jag bättre .
Jag talar lite skotsk galiska .
Känner jag honom ?
Hur vågar du skratta åt mig ?
Bob kom hit , inte sant ?
Jag hör till basebollaget .
Vi hade en mild vinter i fjol .
God morgon .
Pandor är vackra djur .
Vad har fört dig hit ?
De byggde en bro .
Mannen som hon ska gifta sig med är en astronaut .
Lyssna noga !
Låt oss försöka !
Jag arbetade hårt hela gårdagen .
Jag vet var hon är .
Var är utgången ?
Kan någon annan svara ?
John byggde en bokhylla .
Herr White är ungefär i min ålder .
Det här en present till dig .
Gud är en fantasifigur skapad för att få oss att känna oss bättre om vår okunnighet om vår egen existens .
Iberismen är en rörelse för att ena de iberiska folken och nationerna såsom Katalonien , Kastillien , Portugal , Galicien , Baskien , Andalusien ...
Förlåt för att jag stör , men min bil är trasig , skulle du kunna hjälpa mig ?
Var är du nu ?
Varför är en del översättningar gråa ?
Anledningen till trafikolyckan rapporterades av polisen .
Det är säkert att äta fiskarna .
Det är säkert att äta fisken .
Ju mer jag lyssnar på henne , desto mindre gillar jag henne .
Du stödjer planen , eller hur ?
Han är inte för fattig för att köpa en cykel .
Det fortsatte att snöa i fyra dagar .
Du kommer gilla honom så fort du fått chansen att prata med honom .
Han är inte en av oss .
Hon ringde mig flera gånger .
Den här sortens arbete kräver mycket tålamod .
Polisen genomsökte det huset för att vara säkra på att de stulna skorna inte var där .
Doktorn funderar noggrant innan han bestämmer sig för vilken medicin han ska ge .
Pojken hoppar .
Hästen hoppar .
Flickan hoppar .
Hunden hoppar .
Vem läser ?
Två barn sitter på staketet .
Det här är lätt .
Det här är svårt .
Du jobbar för hårt .
Ta det lugnt en stund .
Han tjänar tre gånger så mycket som jag gör .
Jag har lånat en bil .
Jag har lånat ett bord .
Jag har lånat två böcker .
Talar du svenska ?
Ja , lite grand .
Nej , inte alls .
Förstår du mig ?
Nej , jag förstår dig inte .
Var snäll och tala långsamt .
Tack , jag förstår nu .
Var finns det en telefon ?
Finns det en busshållplats här i närheten ?
Ja , där borta .
Kan jag hjälpa dig ?
Kan du säga mig hur man går till amerikanska ambassaden ?
Ingen orsak .
Kan jag få köpa några vykort ?
Hur många vill ni ha ?
En krona och femtio öre .
Var snäll och ge mig en Dagens Nyheter också .
Hur mycket blir det ?
Det blir fyra kronor , tack .
Vi äter lunch .
Vi äter middag .
Vi äter frukost .
Kan jag få se på matsedeln ?
Kan jag få ett par ostsmörgåsar ?
Vad vill ni ha att dricka ?
Kaffe ?
Kan jag få ett glas mjölk ?
Kan jag få ett glas vatt ?
Kan jag få ett glas öl ?
Kan jag få ett glas vin ?
En kopp kaffe , tack .
En kopp te , tack .
Lite smör och bröd .
Det finns en restaurang här .
Det finns en buss här .
Det finns en krona här .
Det finns en telefon här .
Det finns en smörgås här .
Det finns en hållplats här .
Det finns ett vykort där .
Det finns ett glas där .
Det finns ett par där .
Det finns ett hotell där .
Finns det en telefon här ?
Jag talar svenska .
Greta går till ambassaden .
Du ska tala svenska .
Du kan förstå svenska .
En kopp kaffe kostar en krona .
Kostar en kopp kaffe en krona ?
Herr Berg hjälper dig .
Hjälper du fröken Hansson ?
Du vill hjälpa mig .
Jag hjälper dig .
Jag ska hjälpa dig .
Jag kommer till hotellet .
Jag vill komma till hotellet .
Jag vet att jag inte vet .
Jag släppte in katten i mitt rum .
Min pappa är inte hemma just nu .
Jag ringer honom ikväll .
Linda älskar choklad .
Japan är varmt och klibbigt om sommaren .
Hon har gått och lagt sig .
Jag är förkyld .
Gör som du vill .
Hur är han ?
De gick mot porten .
Han satt och läste en bok .
Räck upp handen om du vet svaret .
Jag har blivit ombedd att informera dig om att din far har dött i en olycka .
Vårt lag besegrade motståndaren med 5-4 .
Jag går alltid .
Jag gick och lade mig lite senare än vanligt .
Jag bad henne att vänta ett slag .
Så långt ögat kunde se var marken täckt med snö .
Alla pojkarna sprang iväg .
Vi sprang hela vägen till stationen .
Han pratade väldigt högt .
Där såg han det han hade drömt om .
En student vill träffa dig .
Jag cyklade enhjuling idag .
Jag känner henne inte alls .
Du verkar ha förväxlat mig med min storebror .
Min väckarklocka ringde inte i morse .
Tom kan köra gaffeltruck .
Har du någonsin ätit japansk mat ?
Alla sittplatser var upptagna .
Jag pluggade i kanske två timmar .
Knulla din mamma .
Jag håller inte med dig på den punkten .
" Lita på mig " , sade han .
Hon stannade fem dagar till .
Du klagar alltid .
Kan vi talas vid i enrum ?
Så romantiskt !
Du borde inte äta här .
Jag måste ställa en dum fråga .
Jag är kär i dig .
Han står på scenen .
Jag ser inget !
Bob var inte med på planen .
Har du någonsin varit på Koreahalvön ?
Jag skulle vilja lägga undan mina ägodelar .
Det ser ut att bli regn .
Han verkade trivas med sitt liv och sitt arbete .
Våren är min favoritårstid .
Jag har inget emot att göra hushållssysslorna .
Jag går hellre än att ta bussen .
När man talar om trollen står de i farstun .
När man talar om trollen .
Pojken var så trött att han inte kunde ta ett steg till .
Man kan lära sig många ord genom att läsa .
Vår fotbollsmatch kommer att skjutas upp .
Jag klarar av att försörja min familj .
Den är för liten .
Det är för litet .
Jag måste lämna dig .
Hon blev väldigt arg på barnen .
Det är middagsdags .
Hon antydde att hon kanske skulle studera utomlands .
De är korta och smala .
Skrivbordet är av trä .
Du behöver inte vara rädd .
Han kommer inte att göra dig illa .
Vad kallt det är !
Vad skulle du göra om du såg ett spöke ?
En bläckfisk har tio armar .
Jag var kolugn .
Hon höll just på att skära upp gurkor .
Vilken lång gurka !
Jag har en ärta i min högra näsborre .
Förr trodde man att bara människor kunde använda språk .
Jag åkte till Europa via USA .
Vira en sjal om ditt huvud .
Att simma över sjön tog nästan kol på mig .
Var är Tom född ?
Min far varken röker eller dricker .
Det var snällt av dig att hjälpa mig med läxan .
Ät mer grönsaker .
Var snäll och stäng av teven .
Jag talar spanska med Gud , italienska med kvinnor , franska med män och tyska med min häst .
Sen sjöng jag en dum låt om en myra som försökte brottas med ett tuggummi .
Jag köpte en grön soffa igår , men den gick inte in genom dörren , så jag fick lämna tillbaka den .
Det där måste vara historiens rödaste finne .
Finns det någon som kan hjälpa mig ?
I fjol var april den varmaste månaden .
Apelsiner innehåller mycket C-vitamin .
Mitt skägg växer snabbt .
Han tabbade sig på jobbet och fick sparken .
Om du tror att du kan locka mig med chokladmjölk , så har du fel , för jag är laktosintolerant .
Hon har en ödletatuering på låret .
Trafikljuset slog om till rött .
Peking är större än Rom .
Peking förändras så fort .
Jag såg på när de flådde en människa den dagen .
Bilden är verklighetstrogen .
Jag skriver en uppsats om franska revolutionen .
Får jag också komma ?
Jag är vegetarian .
Gjort är gjort .
Har du gått ner i vikt ?
Hennes röst går mig på nerverna .
Stormen har orsakat fruktansvärda skador .
Jag vet bara inte vad jag ska säga .
Berätta för mig .
Han arbetar hårt året runt .
Trädgårdsmästaren planterade en ros mitt i trädgården .
Jag spelar ofta volleyboll .
Så vitt jag vet håller de alltid sina löften .
Du är röd i ansiktet .
" Det brinner ! " skrek han .
Nästan tre .
Det finns ett parallellt universum i Bermudatriangeln .
All kunskap är inte till godo .
Är Ginza Japans livligaste gata ?
Finns det något bord för två ledigt på fredag ?
Ta fram din plånbok .
Jag har inga pengar på mig .
Hunden har bitit hål på min ärm .
Han är från England , men är väldigt dålig på engelska .
Han är på väg att gå .
Han kunde inte gå längre .
En lång tystnad följde .
Jag är orolig för hennes hälsa .
Får jag låna ditt suddgummi ?
Han erkände sina misstag .
Det var du som föreslog att vi skulle se den filmen .
Vem skrev brevet ?
Ingen annan än du kan göra mig lycklig .
Hur lång är den där bron ?
Soldaten uppgav sitt namn .
Om han ansträngde sig så skulle han lyckas .
Grannhunden skäller alltid .
Mjölken håller i två dagar .
Var snäll och gå till kirurgavdelningen .
Vi bor nära stationen .
Du måste vara jättehungrig nu .
Han har dussintals böcker om Japan .
Hon skyndade ner för trapporna .
Förresten , spelar du fiol ?
Det haglar i regel om sommaren .
Det sade du inte .
Vem är hon ?
Han verkar förakta folk från Kakogawa .
Han tjänar inte mer än femtio dollar i veckan .
Jag åker till Hiroshima tre gånger i månaden .
Har du skor och strumpor ?
Som tur är blev ingen blöt .
Där är Tokyo .
Jag ber om ursäkt om jag har sårat dig .
Jag fryser .
Kan jag stänga fönstret ?
Jag letar efter min nyckel .
Jag säger det hela tiden .
Kan du bevisa det ?
Generalen visade mig vilka kort han hade på handen : spader kung , spader dam och ruter knekt .
Min dröm är fortfarande bara en dröm .
Först trodde jag att han var lärare , men det var han inte .
Jag hoppas att din förkylning går över snart .
Jag ska gå rakt på sak .
Du får sparken .
Han är min bror , inte min far .
Han är lärare .
Vi hoppas på fred .
Jag diskar .
Vi är människor .
Hon målar varje dag , oavsett hur mycket hon har att göra .
Fråga henne vad hon har köpt .
Han skrev ner sina tankar i sin anteckningsbok .
Diamanten värderades till 5 000 dollar .
De här skorna passar perfekt .
Jag är upptagen med maten för tillfället .
Han skrev ner telefonnumret .
Det beror helt på huruvida de kommer att hjälpa oss .
Vi känner till legenden om Robin Hood .
Han är inte här längre .
Man trodde att valar var fiskar .
Tom dömde en konsttävling .
Jag är hans vän och kommer så förbli .
Hon borde ha gjort klart sina läxor .
Spädbarnet log mot mig .
Italiens befolkning är hälften så stor som Japans .
Det här är min fru , Edita .
Mitt hår är längst i klassen .
Han levde inte upp till förväntningarna .
Vi besökte historiskt intressanta platser .
Vad sägs om en kopp kaffe ?
Hon blev påkörd av en bil .
Han är nöjd med sin nya bil .
Hon har många vänner i Hongkong .
Den stackars hunden slets bokstavligen i stycken av lejonet .
Jag pratar inte med dig ; jag pratar med apan .
Vad är klockan ?
Min klocka går fel .
Känner du till någon bra restaurang ?
Jorden är ingen stjärna , utan en planet .
Det kommer inte göra ont .
Min klass består av fyrtio studenter .
Följden blev att hon förlorade jobbet .
Pojkar härmar ofta sina idrottshjältar .
Jag försörjer min familj .
Det tog en månad för min förkylning att gå över .
Sen då ?
Jag avskyr att se djur lida .
Kanske förstår hon senare vad jag menade .
De har en gemensam hobby .
Döm inte andra efter dig själv .
Du måste intressera dig för aktuella händelser .
Håll käften , annars åker du ut .
Förenta nationerna är en internationell organisation .
Jag tycker om att läsa innan jag går och lägger mig .
Det är ingalunda lätt att bemästra ett främmande språk .
Jag tog med mig min kamera .
Sitt inte på den där bänken är du snäll .
Jag skulle vilja följa med , men jag är pank .
Var snäll och ge oss två knivar och fyra gafflar .
Jag är mätt .
Hon ser ut att vara full .
Vi blev stupfulla .
Och slutligen , tolv poäng till Estland !
Kaniner tycker om morötter .
Vill du inte simma idag ?
Den här stolen är väldigt bekväm .
Det är inte lönt att försöka lösa det här problemet .
Det är ingen mening med att försöka lösa det här problemet .
Jag gick inte , utan stannade hemma .
Vem vet inte ?
Jag står inte ut med oljudet längre .
Det är ingen bra bil , men det är en bil .
Vill du ha lite mer sås ?
Golden Gate-bron är gjord av järn .
Hon vann första pris i en matätartävling .
Herregud , jag tror inte det är sant .
Frihet kostar .
Juryn är oenig .
Prata långsammare .
Han såg en hund i närheten av dörren .
Är din mor hemma ?
Pojken tömde tallriken på ett ögonblick .
Jag vill dö med Getter Jaani .
Religion är ett opium för folket .
Hon vill hålla honom på avstånd .
Jag hann precis med sista tåget .
Nu är det lagom , varken för tungt eller för lätt .
Du äcklar mig .
Is smälter i vatten .
Min bror bor i en liten by .
Tre öl och en tequila tack !
Jag tycker att vi ska vänta en halvtimme till .
Strumporna luktar illa .
Då är det dags för din halshuggning .
Har du inga sista ord ?
Han kan inte ens skriva sitt eget namn .
Guld är tyngre än silver .
Hennes far avled i förra veckan .
Jag har inte sett av honom på ett tag .
Han somnade med radion på .
Råttor förökar sig fort .
Den här filmen är sevärd .
Jag skulle vilja hyra en bil .
En bild säger mer än tusen ord .
Var är de andra flickorna ?
Byggnaden totalförstördes i jordskalvet .
Jag tycker om att gå och titta på baseboll .
Hunden grävde en grop .
Hon ville gifta sig omedelbart .
Vi blir tvungna att skjuta upp matchen till nästa söndag .
Han blåste på sina fingrar för att värma dem .
Jag har svårt att tro på det .
Vi måste försvara vårt land till varje pris .
Det här kommer att bli den varmaste sommaren på trettiosex år .
Jag tar det här paraplyet .
Mötet avslutades vid lunchtid .
Kunskap är makt .
En gång i tiden trodde man att människor inte kunde flyga .
Trots att det regnade ställdes matchen inte in .
Vatten , tack .
Skratt smittar av sig .
Men vad vill du ?
Sömnbrist är inte bra för kroppen .
Vi kommer alltid att vara tillsammans .
Hönan har värpt ett ägg .
Han har det bättre än någonsin .
Kan du latin ?
Var är tidningen ?
De lade ut mattan på golvet .
Vad är skillnaden mellan en duva ?
Hon läste hans brev om och om igen .
Jag kan inte böja min högerarm .
Hur smakar den här soppan ?
Varför inte ansöka om jobbet som tolk ?
Vi råkade befinna oss på samma buss .
Hon skämdes för sin obetänksamhet .
Det kanske blir regn snart .
Han höll andan .
I det här fallet tror jag att han har rätt .
Dagarna blir allt längre .
Hon ser fram emot att få träffa honom igen .
Bränt barn skyr elden .
Det går inte att förväxla honom med hans lillebror .
Jag äter inte kött , fisk , skaldjur , fjäderfän eller buljong .
Det ligger en sax på bordet .
Sten , sax , påse .
Du borde gå till tandläkaren .
Vilken spännande match !
Jag skulle vilja ha två kilo äpplen .
Den gamle mannen satte sig ner .
Ja , så vitt jag vet .
Jag har sett fram emot att få träffa dig .
Jag gissade att hon var fyrtio .
Det tar inte särskilt lång tid .
Jag föddes sådan här !
Jag fick en bot på tjugo dollar för olovlig parkering .
Den här boken finns bara tillgänglig i en affär .
Han satte sig på bänken .
Han blåste ut ljuset .
Fysik är mitt favoritämne .
Hennes arm är gipsad .
Ni har rätt .
Nudelsoppan är ganska dyr här .
Jag har inte så mycket pengar med mig .
Problemet är att pojken aldrig gör vad han blir tillsagd att göra .
Jag återvände till Japan .
Tror du verkligen på spöken ?
Det luktar som om någon har rökt här inne .
Vi ses i skolan imorgon .
Bill är på väg till New York .
Jag besöker honom varannan dag .
Jag hör ett konstigt ljud .
Han lever i lyx .
Kom när du vill .
Det finns mer än 4000 språk i världen .
Hawaii har fint väder året runt .
Huset omgavs av en stenmur .
Han är vid hennes sida .
Frågan var omöjlig för oss att besvara .
Vi ska se en utländsk film ikväll .
Kan du inte skilja på fantasi och verklighet ?
Får jag gå på toaletten ?
Han sparkade in bollen i mål .
Mayuko kan cykla .
Han har glasögon .
Jag var irriterad över att hon fortfarande sov .
I Europa startar skolorna i september .
Vad vill du köpa ?
Pandor bor i bambusnår .
Har Bob rätt ?
Tre studenter .
Här är min studentlegitimation .
Du har rätt .
Jag tar en taxi .
Han tvingade sig in i rummet .
Många ryssar krävde ett slut på kriget .
För länge sedan besökte jag Kanada .
Jag somnade .
Förresten , hur många av er för dagbok ?
Jag är i bilen .
Jag är helt säker !
Jag har varit här sedan klockan fem .
Hon är ute efter ett bättre jobb .
Grekiska filosofer värderade demokrati högt .
Kan du säga det en gång till ?
Han gick till affären för att köpa lite apelsiner .
Den här maten luktar ruttet .
Jag är ganska trött idag .
Han använde hennes cykel utan att fråga om lov .
Jag är orolig för honom .
De fångade räven med en fälla .
Hon har ännu fler böcker .
Kortkorta kjolar har blivit omoderna .
Kassören stoppade kundens varor i en påse .
Hennes hår är långt och vackert .
Inte så mycket senap .
Jag stannar här tillsvidare .
Många tror att jag är tokig .
Bara du kan göra detta .
Berätta något om ditt land .
Jag måste bege mig nu .
Hon är väldigt rädd för ormar .
Min mormors sjuksköterska är väldigt snäll .
Min farmors sjuksköterska är väldigt snäll .
Advokaten förklarade den nya lagen för oss .
Vad vill du att jag ska prata om ?
Han höll henne i ärmen .
Jag ringer dig vid sju .
Han beundrade min nya bil .
Kate har tyska som huvudämne .
Tyvärr , jag har ingen aning .
Hjälp mig lyfta paketet .
De såg efter pojken .
Han viftade bort flugorna .
Du får inte formatera den här disketten .
Har man sagt A , får man säga B.
Hon rörde om i kaffet med en sked .
Han är tillbaks om några dagar .
Repet gick av medan vi besteg berget .
Ur vägen , pojk .
Hur länge har du varit utomlands ?
Han är min bror .
Vilka underbara blommor !
Byggnaden uppe på kullen är vår skola .
Det är en present till dig .
Vem som helst kan göra misstag .
De stod på rad .
Katter tycker inte om vatten .
Jag har aldrig ätit mango förut .
Hon var på väg att svimma .
Såg du blicken han gav mig ?
Jag är högerhänt .
Jag hörde dörren stängas .
Jag gillar främmande språk !
Sverige hade chans att ta VM-guldet i ishockey , men förlorade stort i finalkampen i Bratislava .
Storleken har ingen betydelse .
Han skrev ner det för att inte glömma det .
Jag vill dricka mjölk .
Det tog mig tre dagar att läsa den här boken .
Midori åt flest apelsiner .
Han går i tionde klass .
Det var bara ett skämt .
I hur många minuter ska jag koka den här frusna sparrisen ?
Jag har stånd .
Tålmodighet är den vackraste dygden .
Jag vet inte vad han har råkat ut för .
Jag vet inte vad som har hänt med honom .
Hon gav honom en massa pengar .
Håll utkik efter hans senaste film som kommer ut nästa månad .
Tillåt inte dig själv att bli tjock .
Betty är danslärare .
Vilken av de två är tyngst ?
Gå upp för den här trappan .
Hon hjälpte dem med bagaget .
Det tog hela kvällen .
Vad jag vill ha nu är en varm kopp kaffe .
Han deltog i mötet .
Soporna ger ifrån sig en förfärlig stank .
Det var hans eget fel .
Han gräver sin egen grav .
Jag gillar verkligen inte Apple-produkter .
Hennes klänning såg billig ut .
Att flyga drake kan vara farligt .
En dag skulle jag vilja äga en segelbåt .
Jag är trött på att äta på restaurang .
Hans stackars hund lever fortfarande .
Släpp in lite frisk luft .
Efter söndag kommer måndag .
Det här rummet är allt annat än varmt .
Du har inget att vara arg över .
De tackade Gud .
Det finns en sjö öster om byn .
Han var i Frankrike .
Drogens effekter är intensiva men kortvariga .
Mitt hus ligger tio minuters gångväg från stationen .
Det regnade kraftigt hela dagen .
Jag studerar konsthistoria .
Det är rea på pälskappor .
Skulle du vilja spela tennis på söndag ?
Här är mitt kvitto .
Finns det en bensinmack i närheten ?
Det är dags för mig att gå .
Det här skrivbordet som jag köpte igår är väldigt stort .
Han skulle hellre dö än att gå upp tidigt varje morgon .
Han har medlemsprivilegier .
Läraren välkomnade de nya studenterna .
Kan du förklara vad det här är ?
Jag kan inte stänga av duschen .
Kan du kolla det åt mig ?
Det läker av sig själv .
Tvätta händerna innan du äter .
Vilken sorts vin rekommenderar du ?
Vad vet du om honom ?
Tom är en duktig cricketspelare .
Han gick motvilligt för att träffa henne .
Betyder det att du vill göra slut ?
Presidenten har avskaffat slaveriet .
Vem vinner ?
Koka ett ägg .
Jag är inte säker på om det här är rätt .
Hon har äntligen nått Arktis .
Meg köpte en burk tomater .
Glöm henne .
Du får bara prata engelska .
De gjorde en märklig upptäckt .
Om man äter för mycket blir man tjock .
Om du äter för mycket kommer du att bli tjock .
Ann spelar ofta tennis efter skolan .
De här är pojkar och de där är flickor .
Se upp för ficktjuvar .
Hissen verkar vara trasig .
De kan tänka och tala .
Det är regnsäsong .
Problemet med honom är att han är lat .
Är den här platsen upptagen ?
Jag har ryggont .
Jag har ont i ryggen .
Hur ofta äter du fisk ?
Jag har läst ut boken .
Jag behöver en kniv .
Vi använder ätpinnar istället för kniv och gaffel .
Lucy kan inte använda ätpinnar .
Snart är det vår .
Jag drömde om honom .
Jag spelar fiol .
Jag vet inte vad klockan är .
Den här boken är för mig vad Bibeln är för dig .
Det visste jag inte .
Hon köpte en kamera till sin son .
Kastanjer måste kokas i minst femton minuter .
Han rensade gatan på kastanjer .
En ekorre gömde sig bland grenarna .
Kaniner är besläktade med bävrar och ekorrar .
Hún eldar illa .
Det har varit en mycket svår vinter .
Jag heter inte " flicka " heller .
Planet har nyss lyft .
Min far är så att säga en vandrande ordbok .
Jag är Lin .
Du verkar frånvarande .
När kommer du tillbaka ?
Ett år senare föddes Paul .
Hon klappade sin son på axeln .
Varför är de här ?
Inte förrän då fick han reda på sanningen .
Tack , det var allt .
Det var ett misstag från deras sida .
Jag gick en konstkurs i fjol .
Jag kan inte besvara din fråga .
Vi är inte amerikaner .
Hon räckte upp handen för att få bussen att stanna .
Jag vet inte hur man köper en biljett .
Hon hjälpte sin far med trädgårdsarbetet .
Det är femtio kilometer till Paris .
Finns vi ?
Ibland är det svårt att skilja rätt från fel .
Som tur är var vädret bra .
Dags att stiga upp .
Hon såg ledsen ut .
Jag känner inte för att äta någonting idag .
Pandor är väldigt smarta .
Hon kom jävligt sent .
New Yorks gator är väldigt breda .
Han är min typ !
Och varför frågar du ?
Jag vet egentligen inte .
Jag vet inte riktigt .
Vi satt mitt i rummet .
Han kom till New York för att söka jobb .
Vi fick aldrig någon tydlig förklaring på mysteriet .
Du pratar för mycket .
Det här är inte min åsikt , bara min översättning !
Du borde ha besökt Kyoto .
Glöm det .
Det är omöjligt att veta vad som kommer att hända i framtiden .
Var har hon lärt sig italienska ?
Jag ser fram emot att få träffa dig nästa söndag .
Han är välavlönad .
Har du ringt henne än ?
Vi har fem sorters grillspett .
Mitt huvudämne är europeisk medeltidshistoria .
Jag är vänsterhänt .
Alla verkar gilla golf .
Han är antingen full eller tokig .
Vi måste avsluta det här arbetet till varje pris .
Han räknade ut ljusets hastighet .
Lättare sagt än gjort .
Jag frågade vem han var .
Du gamla , du fria , du fjällhöga nord Du tysta , du glädjerika sköna !
Jag hälsar dig , vänaste land uppå jord , Din sol , din himmel , dina ängder gröna , Din sol , din himmel , dina ängder gröna .
Du tronar på minnen från fornstora dar , då ärat ditt namn flög över jorden .
Jag vet att du är och du blir vad du var .
Ja , jag vill leva jag vill dö i Norden , Ja , jag vill leva jag vill dö i Norden .
Han har sålt sin bil , så han tar tåget till kontoret .
De lät mig vänta länge .
Hur vill du ha ditt kaffe ?
Du borde köpa en telefonsvarare .
Jag vet inte vad det här ordet betyder .
En man kom fram till mig och bad om en tändsticka .
Jag vill ha fläkten .
Sysslar du med någon sport ?
De kommer inte förrän imorgon .
Nancy tycker om inomhussporter .
Du måste ta tjuren vid hornen !
Jag behöver en låda i den här storleken .
Deras kontor visade sig ha många kvinnor .
Memorera dikten till nästa vecka .
Det visade sig vara sant .
Jag hittar inte min portfölj .
Det här är det sötaste spädbarnet jag någonsin har sett .
Hunden vill gå ut .
Hon är mörkhyad .
Hanako har glömt sitt paraply igen .
Trots sin sjukdom gick han ofta till jobbet .
Den nuvarande regeringen har många problem .
Huset är målat i vitt .
Han är galen i baseboll .
I morse klarnade det .
Han bar sig illa åt .
De hårda kraven är ett villkor för att Grekland ska få de 60-70 miljarder euro som behövs för att undvika en statskonkurs .
Nu har de tre barn .
En av fördelarna med att bo i en demokrati är att man får säga vad man tycker och tänker .
Presidenten är för närvarande i Miami .
Det är svårt för mig .
Inga stjärnor syntes på himlen .
Jag har ingen aning om hur man spelar golf .
Han berättade sanningen .
Han sade sanningen .
Lugna ner dig .
Lugna ner er .
Vad finns i den här lådan ?
Det där är inte en gul krita .
Hjärnan är bara en komplex maskin .
Jag är nöjd med de här skorna .
Medan han pratade hördes ljudet av ett skott som avlossades .
Medan han pratade hördes ett skott avlossas .
Jag tar ett bad varannan dag .
Jag duschar varannan dag .
Att höra är att lyda .
Pilla inte på såret .
Långa kjolar är på modet .
Du måste inte äta .
Jag är så lycklig !
En fladdermus är lika lite fågel som en råtta .
Var försiktig så att du inte blir förkyld .
Vad gjorde du förra söndagen ?
Han högg ned det där körsbärsträdet .
Här är mitt visitkort .
Du gillar visst inte sashimi ?
Det här är en vän till mig .
Kom du med första tåget ?
Han behöver en stege .
Får jag prova den här ?
Jag har en fruktansvärd tandvärk .
Släpp inte taget .
Din dotter går på droger .
Jag ger mig av nu .
Vart fan ska du ?
Jag hittar inte det jag vill ha .
Det rådde brist på importerad olja .
Men han ville väldigt gärna ha en son .
Han sade till henne att han älskade henne .
Hotellet drivs av hans farbror .
Hotellet drivs av hans morbror .
Han kunde inte förmå sig att skjuta hjorten .
Kan du inte skriva med kulspetspenna ?
Hon svor högt .
Han har setts som Japans svar på Picasso .
Jag har en vän vars far är en känd pianist .
Han bestämde sig för att en gång för alla sluta röka .
Han lämnade boken på bordet .
Magdalena och Ania är goda vänner .
Både Magdalena och Ania är från Polen .
Tímea är en ungrare som bor i Polen .
Det saknas en gaffel .
Vad gjorde du i helgen ?
Hon böjde sig ner .
Jag hade hans namn på tungan , men jag kunde inte komma ihåg det .
Tom samlade på kaffekoppar .
Jag följer inte med .
Hon har känt honom länge .
Hon såg upp mot himlen .
Han låg på rygg .
Det är inte lönt att klaga .
Din högra strumpa är utochinvänd .
Jag hittar inte Tim .
Folk älskar frihet .
De har något gemensamt .
Ät så mycket du vill .
Var har bildats i såret .
Hans fel var avsiktligt .
Vi singlar slant om det .
Jag är skyldig honom 100 yen .
Rökning dödar .
Hon beställde en kopp te .
Jag vill tro att jag vet vad jag pratar om .
Han bestämde sig för den röda bilen .
Jag stannar här till i övermorgon .
Ubåten var tvungen att bryta igenom ett tunt istäcke för att kunna gå upp till ytan .
Sydde du den här för hand ?
Jag växte upp på landet .
Hur dags gick du och lade dig igår ?
Jag tycker bättre om roliga filmer .
Jag tog mig friheten att ringa henne .
Jag kunde inte sova .
Hinner du ?
Hur reagerade hon på nyheten ?
Du då ?
Jag tror det är dags för mig att dra .
Den största skillnaden mellan bandy och innebandy är att bandy spelas på is .
Har du skrivit klart din uppsats ?
Ishockeypucken är inte sfärisk .
Vi drack soju i karaokebaren .
Koreaner tycker inte om koriander .
Finns det ingen annan metod ?
Jag vill komma i kontakt med henne .
Är du ledig i eftermiddag ?
Han ser lite trött ut .
Jag behöver ett jobb .
När fick du konsertbiljetten ?
Du har spillt lite ketchup på din slips .
Ett kilo ketchup motsvarar två kilo tomater .
Soldaterna var utrustade med vapen .
Var kan jag få tag på kartan ?
Visst är det vackert väder ?
Jag vill studera utomlands .
Jag vill plugga utomlands .
Jag tror inte att han kommer .
Studenterna delade in sig i tre grupper .
Jag åt snabbt upp min lunch .
Köpte du den på svarta marknaden ?
Träffade du honom ?
Behöver jag någon medicin ?
Jag känner inga blinda män .
Prinsessan låg och blundade .
Hans bok blev föremål för kritik .
Jag är van vid att jobba hårt .
Vilken frukt tycker du bäst om ?
Ben har också något med saken att göra .
Jag är inte intresserad .
Först till kvarn får först mala .
Stör inte Tom medan han läser .
Länge leve konungen !
Finns det en tvättmaskin i huset ?
Jag bor intill leksaksaffären .
Det är iskallt .
Den här klubben har femtio medlemmar .
Vi turades om att köra .
Alla äpplen som faller till marken äts upp av grisarna .
Hon verkade inte intresserad .
Ställ undan cykeln .
Jag vill att du håller ditt löfte .
Vet du vem som har skrivit den här romanen ?
Vi ska mötas vid sju .
Vi såg många skepp i hamnen .
Olyckor av det här slaget sker ofta .
Hon kanske inte kommer .
Floden är femtio meter vid .
Har du någon legitimation ?
Var är chefen ?
Var snäll mot henne .
Vad kostar den här radion ?
Det tog honom tre månader att lära sig cykla .
Att filosofera är att lära sig dö .
Min hund låtsas ofta sova .
Vi bryr oss inte om vad han gör .
Hans tal var för kort .
Troligt är att inget språk fullständigt saknar lånord .
Du är fortfarande ung .
Vem röstade du på i valet ?
De vägrade låta tågen röra på sig .
Han spelar golf .
Vi hinner med tåget .
Du hinner inte i tid till skolan .
Tror du vi hinner i tid till flygplatsen , Paul ?
Jag behöver skölja munnen .
De är min farfars böcker .
De är min morfars böcker .
Morfar pratar väldigt långsamt .
Farfar pratar väldigt långsamt .
Min farfar hör lite dåligt .
Min morfar hör lite dåligt .
Jag tar hand om min farfar .
Jag tar hand om min morfar .
Hör du fåglarna sjunga ?
De stal min vinflaska !
Han började gråta .
Jag känner mig som en annan person .
Jag tror hon är 40 år .
Vänta , skojar du ?
Varför skulle vi vilja åka till en sådan avlägsen plats ?
Behöver jag opereras ?
Jag lyssnar på musik .
När jag väl öppnade ögonen igen satt Amina och stirrade på mig genom botten av sitt ölglas .
Det var min tur att städa rummet .
Vad heter den här gatan ?
Hunden bet mig i handen .
Grodan och jag turades om att gissa vad det hemliga receptet var .
Har du badat än , Takashi ?
Trottoarerna var blöta efter regnet .
Många vackra blommor blommar på våren .
De flesta slott omges av en vallgrav .
Prata inte strunt .
Jag vill ha pengarna tillbaka .
Hon har en fin docka .
Det värsta med sommaren är värmen .
Det värsta med sommaren är hettan .
Jag är uppe och står igen när mitt ben har läkt .
Han kastade ut mig ur huset .
Jag är ingen morgonmänniska .
Jag hittade ett jobb åt honom .
Japan och Sydkorea är grannländer
Vad heter du ?
Du behöver inte ta av dig skorna .
Hon hade en radio .
Hennes engelska är utmärkt .
Du dödar mig långsamt .
Kommer dag , kommer råd .
I mörkret är alla katter grå .
En liter mjölk innehåller ungefär trettio gram protein .
Jag var ung och jag ville leva .
Jag mådde dåligt .
Ursäkta , vad är klockan ?
Jag har trott på Kylie Minogue sedan 12 juni 1998 .
Talar du turkiska ?
Hon fortsatte prata .
En av oss två måste göra det .
Jag tycker att din engelska har blivit mycket bättre .
Jag har stängt alla sex fönster .
Jag kan inte tacka nog för din vänlighet .
Verklighet och fantasi är svåra att skilja på .
Till min förvåning så hade han en vacker röst .
Denna bok duger .
Den här boken duger .
Det är farligt att bo bredvid en vulkan .
Han tycker om djur .
Min ordbok är mycket användbar .
Det här är den kallaste vintern som vi har haft på trettio år .
Två tredjedelar av eleverna kom till mötet .
Borde jag köpa någonting till honom ?
Det där är poeten som jag träffade i Paris .
Vem skrev det här brevet ?
De är vegetarianer .
Ingenting kan inte existera , för om det gjorde det så skulle det vara någonting .
Man ska inte väcka en sovande orm .
Min åsikt skiljer sig från din .
Han blev tilldelad en ansvarsfull position .
Efter klockan 11 så började gästerna att bege sig av i grupper om två och tre .
Jag protesterade när kyparen försökte ta min tallrik .
De ser honom som en hjälte .
Hur många böcker äger du ?
Dammen har torkat ut .
Gud skapade världen på sex dagar .
Jag har inte tid att göra mina läxor .
På sistone har jag inte haft tid att läsa böcker alls .
De rika är inte alltid lyckliga .
Jag älskar arabiska .
Efter tio minuter så var hon på andra sidan .
Är du okej ?
Detta är en häst .
Många bäckar små blir en stor å .
Är du trött ?
Jag är jättetrött men vill inte gå och lägga mig .
Jag har bara smör i kylskåpet .
Det finns mjölk i kylskåpet .
Finns det nåt att drycka i kylskåpet ?
I morgon ska jag åka till Amerika .
Den här pojken har en stark , sund kropp .
De leker gärna i snön .
I länder som Norge och Finland har de mycket snö på vintern .
Sverige har sitt eget språk .
De kommer från Sverige .
Du kommer från Sverige .
Bron mellan Danmark och Sverige är nästan fem mil lång .
Sveriges befolkning ökar .
Vi tillbringade en utmärkt semester i Sverige .
Jag kommer från Norge .
Bajkalsjön i Ryssland är världens djupaste sjö .
Vladivostok är en stad i Ryssland .
Det här landet heter Ryssland .
Han talar perfekt ryska .
Ryssland blev en andra supermakt .
Den här författaren är rysk .
Moskva är en rysk stad .
Hon talar ryska .
Han talar ryska .
Han kan också tala ryska .
Vi lär oss om antikens Rom och Grekland .
Det var en gång en stor konung som bodde i Grekland .
Min far hade redan varit en gång i Grekland .
Det finns många öar i Grekland .
Turkiet var starkare än Grekland .
Många unga romare åkte till Grekland .
De döpte hunden till Shiro .
Jag ser ett hus .
Träden är gröna .
Det var en gång en fattig man och en rik kvinna .
Det var en gång en grym konung .
Hon läste inte boken .
Han skrev till sina föräldrar .
Talar du hebreiska ?
Det finns ett äpple på bordet .
Jag förstår mig inte på musik .
Får jag äta detta ?
Han tycker att lyssna på radio .
Välkommen !
Tycker du om japansk maten ?
Du kan välja vilken du vill .
Hans hus var litet och gammalt .
Du kom inte till skolan i går .
Jag behöver kompisar .
Om du vill vara fri , försttör då nu din TV .
Jag älskar det occitanska språket .
Vi ska se .
Jag är kines .
Vilken frukt är röd ?
Detta är min vän Tom .
I begynnelsen skapade Gud himmel och jord .
Har man sett på maken !
Se så .
Var är äpplen ?
Nordkoreas tillbakadragne ledare besöker Ryssland för förhandlingar om energi .
Han beskrev i detalj vad som hade hänt .
För tillfället har jag inte nog med pengar .
Jag skrev ner hans namn för att jag inte skulle glöma det .
När Marko kom , sov jag .
Bob har flera böcker i sitt rum .
På min nästa besök tar jag blommar med .
Den här filmen är för barn .
Jag är kvinna .
Ett piano är dyrt .
Hon gav mig de här gamla mynten .
Hon gjorde en kovändning .
Hans tal rörde oss .
Vad är skillnaden på ett piano och en fiol ?
Ett piano brinner längre .
Hej världen !
I dag var havet varmt !
Jag har bröder .
Tom är annorlunda .
Den såg billig ut .
Tycker du om japansk mat ?
Han är trött på mina problem .
Jag kan inte tacka dig nog för det du gjorde för mig .
Jag är lärare .
Det är en fin dag .
Hon är stark .
Det är en sjukdom som inte kan förebyggas .
Tom kom för att be oss om hjälp .
Hon frågade var huset låg .
Min mamma kan inte läsa utan glasögon .
Jag måste göra klart läxan innan middagen .
Herr Yoshida har aldrig brutit ett löfte .
Han sade att han låg sjuk , vilket inte var sant .
Jag skämdes .
" Vad är det som händer i grottan ?
Jag är nyfiken . "
" Jag har ingen aning . "
Mjölk är en vanlig dryck .
Jag går till arbetet varje dag .
Det är allt annat än omöjligt .
Jag är japan , men du är amerikan .
Det är skönt att stiga upp tidigt .
Det var snudd på otänkbart att pojken skulle stjäla .
Han gick ut trots ösregnet .
Tom kunde knappt förstå vad Mary sade .
Tom är granne till Mary .
Man måste dra gränsen någonstans .
Han är lång och stilig .
Allt du behöver göra är att trycka på knappen .
Jag spelade tennis med min bror .
Är det din egen idé ?
Var snäll mot andra .
Tro på dig själv .
Papegojan är död .
Guld är mycket tyngre än vatten .
Det är en harpa .
Nunnorna sjunger .
Din önskan har gått i uppfyllelse .
Jag promenerar till jobbet varje dag .
Utsikten är fantastisk .
Jag är i San Diego och ni bara måste komma och hälsa på mig !
På inrådan av sina astronomer bestämde sig Alexander den store för att inte attackera Egypten och for till Indien istället .
Vad kämpar du för ?
Dags att sticka .
Min syster tycker om Ultraman .
Tom öppnade dörren för Mary .
Det är en gammal kvinnas röst .
Jag blödde näsblod idag .
Det är Babas röst .
Jag tappade bort min väska på väg till skolan .
Jag vill inte gifta mig .
Det var inget sammanträffande .
Detta är reglerna .
För att dölja det faktum att hon var en princessa förklädde hon sig till en pojke och flydde från slottet .
Jag har aldrig träffat dig i verkligheten .
Du är trygg här med mig .
Jag med .
Det kan jag inte utesluta .
Det är roligt att spela baseball .
Mina föräldrar är väldigt stränga .
Låter det bekant ?
Jag har fått nog .
Skitsamma .
Ge mig dina tankar .
Jag har stämt träff med honom klockan tolv .
Alkohol löser inga problem , men det gör inte mjölk heller .
Han tvättar bilen .
Jag presenterade mig på mötet .
De betedde sig underligt .
Jag blev blöt ända in på skinnet .
Följ efter mig !
Jag pratade med min farbror i telefon .
Jag pratade med min morbror i telefon .
Det är svårt att skilja sanning från lögn .
Bill lyckades bli godkänd på provet .
Hon såg fram emot att gå på bio med honom .
På grund av några oundvikliga omständigheter i sommar kan jag inte bo i min semesterstuga .
Gnugga fläcken med vinäger .
De har tolv barn .
Tyvärr dog hon ung .
Hon tycker om rysk pop .
Hon var försiktig med att inte slå sönder glasen .
Följ den här gatan i ungefär fem minuter .
Tom kan komma på vår fest i morgon .
Tom berättade för Mary om John .
Tom tar en promenad varje eftermiddag .
Det stod i tidningen att ännu ett krig har brutit ut i Afrika .
Jag har fått nog !
Jag har varit död förr , och det var inte så illa .
Det låter som en bra idé .
Han stiger upp klockan sju .
Hon har satt sitt hus till försäljning .
Det ligger affärer längs gatan .
Var snäll och dela ut korten .
Jag skulle inte vilja vara i hennes skor .
Jag tänkte ringa honom , men jag kom på bättre tankar .
Detsamma gäller Japan .
Jag har massor av kameror .
Vad är de gjorda av ?
Jag har bestämt mig för att gå i pension .
Tåget avgår om tio minuter .
Du borde inte gå ut i den här kylan .
Jag är rädd för bussen .
De här kängorna tillhör henne .
Tom tror inte att detta är någon tillfällighet .
Hon måste hjälpa honom .
Inget är omöjligt för Gud .
Tappa inte den där koppen .
Hon har en väldigt prydlig handstil .
Jag vet inte vad rätt svar är .
Jag hatar alla slags insekter .
Du förstör alltid allting .
Hennes söner har åkt till Tokyo .
Hon rådde honom att ta medicinen .
Tom och Mary vaknade tidigt för att se årets första soluppgång .
Hur länge har det snöat ?
Han besökte ett barnhem i Texas .
Du måste sluta ljuga för dig själv .
Den här skolan grundades år 1970 .
De talar spanska i Mexiko .
Nej , jag gick ut .
Du får skriva på vilket språk du vill .
På Tatoeba är alla språk likvärdiga .
Allt är Toms fel .
Du borde inte döma folk efter utseendet .
Man ska inte döma folk efter utseendet .
Vad oroar du dig för ?
Explosionen skakade hela byggnaden .
Jag kunde inte föreställa mig att jag skulle känna såhär för dig .
Vi har diskuterat det här problemet nyligen .
Det här är löjligt !
För Guds skull .
Min dator har hängt sig .
Jar har ett hus i bergen .
Det kommer att ta några dagar att gå in de här skorna .
Trots alla hennes brister gillar jag henne .
Hon kommer aldrig i tid .
Pojken gjorde sig lustig över flickan .
Den här stenen är dubbelt så tung som den där .
Det är något fel på min bil .
Tom bestämde sig för att säga upp sig .
Till slutet av veckan .
Meg ringde efter dig medan du var borta .
Han är grov till sättet .
Tom verkar sova .
När det slutar regna ska vi ta en promenad .
Tom bad Mary hålla ett tal .
En morgon såg han en söt flicka .
Han såg ut som om han vore sjuk .
Hon är på intet vis självisk .
Jag har aldrig blivit kär i någon tjej .
Hon lyckades inte övertala honom till att hålla tal .
Han förblev obesegrad under hela sin karriär .
Du passar bra i kort hår .
Jag fick reda på var hon var .
Har du redan bokat våra platser på flygplanet ?
Jag vill lära mig standardengelska .
Jag tror på hennes berättelse .
Jag läste just ut Svindlande höjder .
Många använder uttagsautomater för att ta ut pengar .
Jag borde ha vetat bättre än att ringa honom .
Tom somnade till slut .
Gick du i skolan idag ?
Han har cancer .
Vilken vacker fågel det är !
Jag har inte tid för dig .
Jag vet att hon har varit upptagen .
Jag har inte tid för er .
Jag skulle vilja att du betalar i förskott .
Den ekonomiska situationen är inte bra just nu .
Den här roboten gör vad jag än säger .
Det är till stor hjälp när jag är för trött för att göra någonting .
Inte alltför troligt , va ?
Den här boken är tung .
Det ska snöa idag .
Han jobbade hårt för att försörja sin familj .
Jag har ont i fötterna .
Hon frågade honom varför han grät .
Min far dog i cancer .
Vi skyndade oss till tågstationen .
Staden grundades år 573 .
Peter är mycket lång .
Han liknar sin far .
Jag träffade honom igår .
Katten sov på bordet .
Han säger att han älskar blommorna .
Hon säger att hon älskar blommorna .
Äter man inte dör man .
Min bror anländer imorgon bitti .
Vi planerar en resa till New York .
Hon är långt ifrån dum .
Hans bil liknar min .
Enligt väderprognosen ska det snöa i morgon .
Den här boken är lika intressant som den där .
Om jag var rik , så skulle jag köpa ett skönt hus .
Han satt på sängen .
Jag försöker lösa det här problemet .
Hur lång är du ?
Toaletten ligger på övervåningen .
Vi har känt varandra i många år .
Huset är i brand .
Igår var det fredag och i övermorgon är det måndag .
Han är stolt över att vara musiker .
Bill talar lite japanska .
Det gemensamma språket bland många asiater är engelska .
De flesta japaner dricker kranvatten .
Skjut inte budbäraren .
Jag beklagar detta missförstånd .
Jag är redo .
Den här kameran är billig .
Jag försökte öppna dörren och dörrhandtaget lossnade .
Han har skrivit många böcker om Kina .
Min son tror på jultomten .
Vad är det här ?
Det här är en stol .
Var hittade du nyckeln ?
Hjälp mig !
Jag kan bo i gästrummet .
Igår eftermiddag skrev jag ett brev .
Bron förbinder de två städerna .
Jag åt med min lillebror .
Han hade massor att göra .
Följer du med mig till affären ?
Vi hade väldigt kul .
Alister dödade Barbare .
Den här bilen drivs av alkohol .
Jag är inte så förtjust i grönt te .
Ställ den var som helst .
Jag lagade kvällsmat .
Det kommer att kosta minst fem dollar .
Jag är typen som skyr risker som pesten .
Vi spelade baseball .
Han är medveten om faran .
Är hon trevlig ?
Jag kom hit tillsammans med mina vänner .
Varje person betalade tusen dollar .
" Är hon ung ? "
" Ja , det är hon . "
Tusentals utlänningar besöker Japan varje år .
Det här är min katt .
Hunden följde efter honom vart han än gick .
Julen närmar sig .
Jag är fortfarande arg på henne .
Hon drömde om vilda jaguarer .
Var god och fyll i detta formulär först .
Tom tror att Mary fattade rätt beslut .
Du borde inte gå ut .
Det kommer att ta tre månader för vår nya skolbyggnad att bli färdig .
Jag oroar mig över hans hälsa .
Jag studerar koreanska .
Fotnoterna finns längst ner på sidan .
Välkommen till mitt liv .
Han dricker för mycket .
Se dig omkring .
Du är anhållen .
Har du pengarna ?
Jag har aldrig varit i Argentina .
Vilken är din favoritsnabbmatsrestaurang ?
Jag är finsk , men jag talar svenska också .
Han hade snö upp till knäna .
Du har bara en chans att svara rätt .
Gör vad du vill .
Det är första min far skrev .
Det trodde jag aldrig om dig .
Vi har ett väldigt allvarligt problem .
Män vet inget om kvinnor .
Det är en papegoja i fågelburen .
Vi kysstes .
Jag tycker om att mata duvorna .
Har du lite bröd ?
Jag ska mata duvorna .
Vi hade en överenskommelse .
Du bröt den .
Minns du den gången vi åkte till Paris ?
Matade du papegojorna ?
Vad är ditt namn ?
Du måste ha blandat ihop mig med någon annan .
Vi har två barn .
Sluta klaga och gör som du blivit tillsagd .
Ta en karta med dig ifall du skulle gå vilse .
Det nuvarande lösenordet är " eosdigital " .
Jag letar efter mina nycklar .
Tom gjorde klart läxan innan kvällsmaten .
Varsågod och sitt ner .
Hunden blöder .
Varför gör du så mot mig ?
Det här är första gången jag skriver ett brev på spanska .
Min bror är lärare .
Trots att jag har läst engelska 6 år i skolan talar jag det inte bra .
Tom är verkligen ledsen .
Han talar lite engelska .
Hur var det ?
Flickan dricker te .
Kommer han hem klockan sex ?
Vilken är nästa station ?
Han låtsas vara döv .
Var hälsad , gillesbroder .
Du är fin i håret .
Skaffa dig ett liv .
Jag hatar dig .
Må balroger äta dig .
En diskret hyllning till olycksoffren hölls igår .
Är det etiskt att ge honom intervjufrågorna i förväg ?
Ett land utan horhus är inget land .
Det finns inga droger här .
Jag gillar utmaningar .
Snabbmat kan vara beroendeframkallande .
Jag har inte tid att laga mat .
Jag vill inte laga mat .
Han hade ont i huvudet .
Det här monumentet restes i februari 1985 .
Låt oss inte tänka så .
Tom sa att han trodde att Mary fortfarande bodde hos sina föräldrar .
Jag skulle vilja åka till Frankrike någon gång .
Han förnekade den uppgiften .
Jag heter Wang Jiaming .
Jag böjer mig inte en millimeter i den här frågan .
Mor stannade i bilen medan far handlade .
Mamma stannade i bilen medan pappa handlade .
Jag kommer inte på hans namn just nu .
Jag ångrar att jag åt ostronen .
Hon såg till att resenären hade mat och kläder .
Hon bar babyn på ryggen .
Vad gör du idag ?
Han steg på tåget .
Hon betalade sju procents ränta på lånet .
Hon har en stuga vid havet .
Det jag inte vill förlora är kärlek .
Filosofi är egentligen hemlängtan ; Längtan att vara hemma överallt .
Fienden kastade in nya styrkor i slaget .
Ju mer vi har desto mer vill vi ha .
Jag hade en besvärlig tid .
Jag hade det besvärligt .
En hund skäller .
Det är skräp .
Släng det !
Om jag visste hennes namn och adress kunde jag skriva till henne .
Det här börjar bli svårt .
Bill hatar att hans far röker mycket .
Min pappa är starkare än din .
Tom gav inte upp .
Det är min bok .
Många människor dödades i kriget .
Hon spelade piano tillräckligt bra .
Han har problem .
John spelade gitarr och hans vänner sjöng .
Jag är dubbelt så gammal som du .
Slåss som en man !
Det här är en rökfri kupé .
Han borde ha varit färdigt nu .
Att förlora min dotter har berövat mig livsglädjen .
Du är en ängel som handlar åt mig .
Han hatar att bli tillsagd att skynda sig .
Så vitt jag vet är han inte lat .
Jag ogillar att vara ensam .
Det blev oavgjort .
Jag uppskattar vår vänskap mycket .
Det är knappast värt att bry sig om honom .
Tåget avgick i tid .
Vem vikarierar för Tom medan han är borta ?
Jag är mycket glad att lära känna er .
Eftersom han ljög straffades han .
Jag föredrar att åka tåg framför att flyga .
Hon har vackra ögon .
Valet låg mycket nära .
Vad gör den här stolen här ?
Tom bär alltid en karta och kompass i sin väska .
Det var en så kraftfull explosion att taket flög av .
Det här svärdet är i gott skick .
Många unga i Japan äter bröd till frukost .
Är vädret fint ?
Mötet varade till 5 .
Vet du varför han skolkade idag ?
Vet du anledningen till att han skolkade idag ?
Hon är utom sig av glädje .
Vad sägs om att stanna ?
Jag visste att jag var tvungen att berätta sanningen för honom , men jag kunde inte förmå mig till det .
Du frågar fel person .
Jag ringer min man .
Jag gillar att gå en tur i parken .
Biljetterna är slutsålda .
Är det nyttigt för dig att äta fisk ?
Han bad om min hjälp .
Han kallades att vittna .
Allt du behöver göra är att vänta och se .
Barnet slutade gråta .
Jag tänker på dig hela tiden .
Vår engelsklärare är både sträng och snäll .
Han är inte vad han utger sig för .
Månen är mycket vacker i kväll .
Jag gör det om du stöttar mig .
Medicinen var hennes sista utväg .
Hur är den nya ledaren ?
Vi väntar främmande i kväll .
Du borde rensa ogräset .
Jag glömde mina bilnycklar .
Till jul har vi känt varandra i tre år
Den ena talar engelska , den andra japanska .
Han var van att flyga ensam och hade i sin fantasi flugit rutten många gånger .
Ge inte upp halvvägs .
Är det utegångsförbud ?
Han föll aldrig för frestelsen .
Denna salen tar 2000 personer .
Jämför de båda noggrant , så ska du se skillnaden .
Jag föreslår honom till ordförande oavsett om du är för det eller inte .
När det regnar såhär får vi aldrig en chans att gå !
Tom satte sig i förarsätet och körde iväg .
Jag är inte ett dugg trött .
Han är bara en vanlig kontorsråtta .
Äpplena han skickade mig var utsökta .
Jag vet var han bor .
Men det är en hemlighet .
Det är svårt för en nybörjare att uppskatta vindsurfing .
När han log , såg barnen hans långa gråa tänder .
Underskottet har minskat lite i taget .
Jag gick inte på grund av sjukdom .
Några är dyra medan andra är väldigt billiga .
Visst är han ung , men han är mycket pålitlig .
Vi kunde inte godta hans berättelse .
Städa golvet med den här moppen , tack .
Hon är kvart över nio .
Det var varmt , och fuktigt till yttermera visso .
Det var varmt och dessutom fuktigt .
Vi såg inga flickor i gruppen .
Vilken föredrar du ?
Den här eller den där ?
Toms nya skjorta krympte i tvätten så nu passar den inte .
Polisen lyckades hitta brottslingen .
Du påminner om en pojke som jag kände .
Hon varnade barnen för att leka på gatan .
Hon har en bild .
Till hans förvåning stannade tåget till kort .
Det finns en park i centrum .
Få saker ger oss så mycket nöje som musik .
Inte en människa syntes till i byn .
Tom slutade röka .
De krävde stränga straff för de södra rebellerna .
Jag yrkar att vi godkänner förslaget och att åtgärder vidtas så fort som möjligt .
Ser du efter barnen medan jag är ute ?
Oddsen för att Reds vinner är 2 mot 1 .
Du har ett meddelande här .
Om någon är politiker är det han .
Om inte människan tar hand om miljön kanske miljön eliminerar mänskligheten .
Tom är ute .
Spring fort , annars kommer du för sent till skolan !
Att äta en klyfta vitlök varje dag , är det nyttigt för dig ?
Han vann matchen tack vare sin starka vilja .
Det är viktigt att följa en sträng diet .
Det är inte söndag varje dag .
Han är på väg och kommer att anlända i sinom tid .
Min far besökte min farbror på sjukhuset .
Aldrig hade jag sett en sådan fridfull syn .
Han var intresserad av Orientens mysterium .
Jag talar japanska väl .
Jag hoppas du har kul .
Tom har något i sin hand .
Han tappade kontrollen över bilen i kurvan .
Jag vill be dig om en tjänst .
En efter en reste sig och gick .
Om det regnar kommer han inte .
Jag har lagat radion åt honom .
Det är risk att du blir en rejäl karl .
Du måste städa ditt rum .
Vi lyssnar med öronen .
Den här whiskyn är för stark .
Vilket märke gillar du ?
Hon har en del egna pengar .
Jag undrar vem som satte igång det där ryktet .
Hon har inte mindre än tolv barn .
Det finns inget annat att göra än att vänta på att platserna blir lediga .
Var får jag tag på böcker ?
Som pojke brukade jag ligga på gräset och titta på de vita molnen .
Jag gillar att ha mycket att göra .
Vi tillbringade en natt i en fjällstuga .
Det finns regler att följa .
Hans sätt var mycket impopulärt .
Min far lagade en trasig stol .
Den långa resan förvärrade hennes skada .
Tom vet inte vad han ska beställa .
Han är bara en flyktigt bekant .
Den andra delen av boken utspelar sig i England .
Fast att vi väntade till tio dök Bill aldrig upp .
Var snäll och vänta en stund medan jag gör klart ditt kvitto .
Bob har många böcker på sitt rum .
Egentligen inte .
Skriver de ett brev ?
Den misstänkte ljög för polisassistenten .
Han såg ut som om inget hade hänt .
Både pojkar och flickor borde studera hemkunskap .
Nyhetsförmedlaren betonar matkrisen för mycket .
Peka inte på andra .
Trots kylan gick vi ut .
Hur kan jag åka buss till sjukhuset ?
Eftersom varorna Ni debiterat oss inte var perfekta kommer vi inte att betala räkningen .
Tjuvar bröt sig in i mitt hus i går kväll .
Det är fritt för fantasin .
Jag behöver den i morgon .
Efter måltiden frågade jag efter räkningen .
Filmen var intressant , precis som jag hade förväntat mig .
Signalen blev grön .
Tom gjorde många misstag .
Han sa ingenting medan jag talade .
Hur länge tänker du stanna här ?
Kom in och sitt ner , är du snäll .
Hon hörde honom sjunga .
Jag har blivit bättre .
Vänta en stund .
Han är angelägen att åka dit .
Jag förstår inte vad du pratar om .
Ingen är för gammal för att lära sig .
Jag undrar varför hon inte berättade om det för honom .
Jag såg på när den röda solen gick ner i väst .
Jag blev tvungen att vänta i tjugo minuter på nästa bus .
Ah , föraren är galen .
Jag kan inte komma på något annat sätt att få honom att acceptera vårt förslag .
Människan som slutar lära sig är så gott som död .
Jag är inte för trött .
Jag är inte på väg någonstans .
Sjön hade frusit till , så vi gick över isen .
Ingen sprang före honom .
Hennes storasyster gifte sig förra månaden .
Han förklarade varför experimentet misslyckades .
Snälla , förlåt mig .
Du kommer att få stå till svars för detta , Ibragim !
John bryr sig inte ett dugg om sina kläder .
Överallt hon kommer är hon uppskattad .
Det där är en bit paj .
Pojken som står vid dörren är min bror .
Tom har inget lokalsinne .
Tom verkar inte vilja sänka priset .
Vi har mycket snö vintertid .
Poängen är huruvida hon kommer att läsa brevet eller ej .
Så du och Hanna planerar att gifta er ?
Jag skulle vilja ha en flaska hostmedicin .
Han är inte sig själv idag .
Jag upprepade vad han sa ord för ord .
Jag gillar sommaren bäst .
Han tycker mycket om musik .
Kumi talade inte om sin klubb .
Han stod på golvet .
Den sjuke ligger i sängen .
Var har du sett de här kvinnorna ?
Du vet inte vem jag är .
Båda vägarna leder till stationen .
Hon gick tjugo mil om dagen .
USA exporterar vete till hela världen .
Hans gamla katt lever fortfarande .
På Esperanto slutar substantiv på " o " .
Plural bildas genom att tillfoga " j " .
På julen äter man gåsstek , rödkål och dumplings .
Jag kände igen henne vid första ögonkastet .
Ingen är perfekt .
Den här stolen är gjord av plast .
Jägaren sköt på fågeln .
Antalet européer som besöker Thailand varje år , är mycket stort .
Fåglar flyger .
Hur gammal är den här hunden ?
Vad läser du ?
Jag har letat efter Andy .
Vet du var han är ?
Vet du hur många människor som dör av svält i världen per år ?
Din mor måste ha varit vacker som ung .
Jag gillar att resa .
Öppna aldrig dörren på en bil i farten .
Ken och Meg är båda två mina vänner .
Som ett sätt att fördriva tiden på en av sina långa resor , bildade Christoffer Columbus en gång en mening med oändligt antal ord .
Vi betraktade honom som ett geni .
Det är emot mina principer .
Jag kommer att ringa för att få det bekräftat .
Esperanto skrivs fonetiskt med hjälp av ett alfabet om 28 bokstäver .
Det är ingen risk för regn idag .
Hon är varken i köket eller i vardagsrummet .
Jag äter en gurka .
Väck det inte .
De här tre vackra flickorna är allihopa mina systerdöttrar .
De här tre vackra flickorna är allihopa mina brorsdöttrar .
Jag tycker mycket om honom , inte för att han är hövlig utan för att han är ärlig .
Prata du på , jag gör som jag vill .
Jag blev uppkallad efter min farbror .
Jag blev uppkallad efter min morbror .
Vem äger den här bilen ?
Fåglarna lägger ägg .
Hur många bokstäver finns det i alfabetet ?
Jag äter kvällsmat kvart över sju .
Jag är alltid stolt över min familj .
Öppna era ögon .
Du beklagar alltid dig alltid över din man .
Då och då studerar jag esperanto .
Från tid till annan studerar jag esperanto .
Hennes flicknamn är Pupkina .
Han är ministern som ansvarar för miljöskyddet .
Det är länge sedan jag såg honom .
Jag behöver hitta ett deltidsjobb .
Du sa att du hade en vacker bak .
Var det bara vilseledande reklam ?
Vänta till trafikljuset slår om till grönt .
Med dig är det sommar året om .
En fet vit katt satt på en mur och betraktade dem med sömniga ögon .
Det skulle ta mig för lång tid att förklara för dig varför det inte kommer att fungera .
Hon har erfarenhet av att ta hand om barn .
Mitt språk är inte med i listan !
Lås dörren !
Fåglar sjunger tidigt på morgonen .
Vindruvorna är så sura att jag inte kan äta dem .
Kan man hitta en telefon i närheten ?
Han är skyldig till stöld .
Var snäll och väck mig klockan sex i morgon bitti .
Strutsar kan inte flyga .
Hur säger man " adjö " på tyska ?
Du ska stanna här till klockan fem .
Jag är riktigt oroad över din framtid .
Varför kommer du så tidigt ?
Tom vet verkligen inte vad han ska göra .
Jag ber om ursäkt för det sena svaret .
Importen av brittiska varor ökade .
Vår plan kommer att fungera bra .
Ett bra vin behöver inte annonseras .
Miljoner vilda djur lever i Alaska .
Hon är pigg på att sticka utomlands .
Reta inte honom bara för att han inte kan skriva sitt namn .
Mor går till sjukhuset på morgonen .
Det är bäst att du inte väntar längre .
I svåra sorgfyllda tider , låt oss då göra något för andra .
Hon är väldigt duktig på att imitera sin lärare .
Sex blev inbjudna , inklusive pojken .
Tom missade chansen att åka till Boston med Mary .
Tom låtsades inte förstå vad Mary sa .
När han åker till Europa kommer han att besöka många museer .
Vem är flickan som står där borta ?
Killen var så barnslig att han inte kunde motstå frestelsen .
Tom samlade ihop alla sina saker .
Jag har förlorat min PIN-kod !
Det går inte att säga hur långt vetenskapen kan ha nått till år 2100 .
Vad i hela världen står på ?
Tar du mig för fyrtio ?
Du missar rejält !
Jag sätter in tiotusen yen varje månad .
Jag sätter in tiotusen yen på banken varje månad .
Ursäkta , kan du förklara vägen till stationen ?
Tom är van att ta snabba beslut .
Han åker om tre dagar .
Han är tillbaka om tio minuter .
Vid hemkomsten upptäckte jag inbrottet .
Vem talar ?
Jag gillar inte modern jazz .
Vi letar efter en nedgrävd skatt .
Vi har en begränsad budget .
Vill du beställa någonting mer ?
Jag är säker på att du lyckas .
Vad krävs för att man ska få lite hjälp ?
Sluta att bita på naglarna .
Det var ett förskräckligt väder .
Han tjänstgjorde utan allvarligare anmärkningar till han uppnådde pension .
Det är Marys tur att diska .
Jag lyckas inte stänga duschen .
Kan du kolla på det åt mig ?
Zürich betraktas som en större finansiell knutpunkt .
Männen gick för att jaga lejon .
Vattnet är rent .
Miljoner människor förstår interlingua vid första ögonkastet .
Dricker du kaffe ?
Gårdagen är historia .
Morgondagen är ett mysterium .
Dagen idag är en gåva .
Det är därför den kallas för nuet .
En dröm är hela livet , själva drömmen drömmer vi .
God jul !
I min värld är alla en ponny , som äter regnbågar och bajsar fjärilar .
En katt har två öron .
Det finns inget ont som inte har något gott med sig .
Barn borde vara nyfikna .
Lätt gånget lätt förgånget .
Som man bäddar , får man ligga .
När PC-fel saktar ner dig , vad kan du göra ?
Många var gråtfärdiga när påven dog .
43-åriga kvinna misstänks ha skjutit ihjäl sin make .
Hovar skrapar i den höstfuktiga ängsmarken .
Jakten på låtsasräven börjar .
Mustasch som ser ut som ett cykelstyre eller bara moppefjun .
Det är bara att välja en överläppsprydnad och testa vad den utstrålar - elegans , töntighet , makt , sexighet eller bara mysfarbror .
Skämtet såg inte ut att falla i god jord hos Sarkozy .
" Tack . "
" Varsågod . "
Kvinnan fastnade på något sätt mellan sin egen bildörr och något annat på uppfarten .
Grekland avblåser folkomröstningen .
Att se regissören Craig Brewers nya tappning av ungdomsklassikern är lite som att återse en gammal förälskelse .
Snubbelhumorn som lärde Hergé sig av stumfilmen .
Ärkeskurken Rastapopolous är en affärsman som inte drömmer om världsherravälde , utan bara om pengar .
När en katt ligger och sover i ett rum finns det inte mycket mer för en inredare att göra där .
Sex får låg döda eller svårt sargade .
Varg eller lo ?
Nej , människa och hund eller möjligen flera hundar hade gått lös på fåren i hagen .
Finansministern , med sin väl tilltagna rondör , tvingades i tisdags uppsöka sjukhus efter att ha fått problem med magen .
Det är ett djupt obehagligt uttalande .
Inte är vi väl så fega , vi som valt att bli idrottsledare att vi inte vågar kritisera varandra , rensa ut rötäggen ?
Premiärministern måsta samsas med andra .
I natt avgjordes regeringens öde .
Hon tål inte ljus , inte ens skenet från en mobiltelefon .
Jag har hållit mitt artisteri lite i skymundan för min familj .
Jag har velat särskilja mig från dem .
Hans karriär rivstartar .
Hon höll på att städa lägenheten .
Visserligen hann inte Chauser klart med hela Canterbury Tales men man räknar ändå den som en av senmedeltidens stora verk .
Köttbullar skulle vara lagom stora , lagom runda och lagom bruna , säger Emils mor .
Han kunde lära sig utan instruktioner .
Städerskan trodde att hon bara gjorde sitt jobb - i själva verket förstörde hon ett modernt konstverk värt miljoner .
Nu brottas museet med hur det ska hantera krisen .
Barnet föddes helt friskt .
Vi vet att han är en modig man .
Man gör leksaker i den här fabriken .
Jag önskar jag kunde köpa det där huset billigt .
Stor förvirring blandat med ilska följde på beskedet från Swedbank nu på eftermiddagen att banken ska göra sig av med 600 anställda .
Herr Smith gläder sig över sin sons framgång .
" Risk för nattfrost på låglänta marker " , sade man i väderrapporten .
En tidigare anställd på ett äldreboende i Staffanstorp döms till villkorlig dom och 10 000 kronor i skadestånd för att ha förskingrat en boendes pengar .
Barn har rätt till en giftfri vardag .
Knep kan ge dig pengar på kontot .
Barn dricker mer vatten , äter mer mat och andas mer luft per kilogram kroppsvikt än vuxna .
Ficktjuven var ovanligt skicklig .
Inte ens en polis på spaningsuppdrag märkte att han blev bestulen på sin Iphone av honom .
Efter avslutat samtal sä ­ ­ ger han vänligt adjö och önskar mig en trevlig kväll .
Nu behöver man vinterdäck .
Det är lätt att glömma att mikrofonen är påslagen .
Det var ett pinsamt fiasko för Rick .
Presidentkandidaten fick hjärnsläpp .
Rysk rymdsond kan krascha .
Experter fruktar giftregn mot jorden .
Det måste du se för att tro på .
Katten var inte längre lika snabb i benen , och en dag hann räven ifatt .
Det var ett pinsamt fiasko .
Gubben var 99 år och fyra månader gammal när han blev bostadslös .
Dessutom saknade han sin katt .
Han vaknade upp till sin hundraårsdag , djupt besviken .
Döda havet lever .
Det lockar turister från världens alla hörn .
Lunds universitet har haft ett problem – för mycket pengar .
Nu har man lyckats sätta sprätt på slantarna .
13-åring krockade föräldrarnas bil .
En svårt hjärtsjuk äldre kvinna återfanns medtagen men vid liv .
Behovet av reformer i Italien är enormt .
Fåren föddes i våren .
Jag hoppas han får ett straff .
Vårdföretag ska inte kunna tysta personalen .
Åter nås vi av nedslående rapporter om missförhållanden i välfärdsverksamheter .
Polisen bluffade om gripna klottrare .
Jag har glömt mina glasögon .
Var har du gömt julklappen ?
” Tekniken är inget hot mot svenska språket ” , säger språkkonsulten Anna Antonsson .
Många tror att unga blir sämre på att läsa och skriva men utvecklingen kan i stället betyda att de får en högre skriftspråklig kompetens .
Flaggor väcker känslor .
Det finns vissa länder där jobchanser för bödlar har tyvärr inte försämrats mycket i de senaste åren .
Det började långsamt , smygande .
Hans hår var kortklippt och han var slätrakad .
Ibland får man bli någon som man tidigare inte var .
Var det inte Kafka som skrev att en bok måste bli yxan för det frusna havet inom oss ?
Han hälsade henne med ett brett leende .
Alzheimers sjukdom börjar långsamt smygande .
En barnkör från grannsocknen sjöng några smöriga låtar .
Nu ska vi ha kalas !
Man kan förändras som människa , men om man byter ut alla sina bästa egenskaper mot nya , så utmanar man ödet .
Det var ett misstag hon brukade undvika med otrolig koncentration .
Tålamodet med Assad är slut .
Det är en film som alla föräldrar borde se .
Det gäller bara att snabbt öppna nya behovslådor och så vips , så måste man ha något nytt .
Trollis försvan spårlöst i vimmlet .
Tomas , 62 , cyklade från surströmmingskalaset .
Katter som springer lösa ute lever farligt .
När den fuktiga vägbanan frös till is bäddade det för blixthalka i länet .
Trädet är ruttet och stendött och kan falla när som helst .
Det rådde god stämning bland de 30 till 40 demonstranter som har samlats .
En riktig cider för mig ska ha en doft av mogna äpplen med frisk äppelsyra och en viss skalbeska – torr med toner av fruktsötma .
Familjen gick vilse i majslabyrint .
Han fick ett hotbrev .
Jag är idel öron .
Jag kan inte komma på någon bra ursäkt till varför jag är sen till tandläkaren .
Kan du simma lika snabbt som honom ?
Han är inte en läkare .
Åh nej !
Mitt hus brinner !
Det var en ny bok .
Vems bok är det ?
Lägg inte plånboken på elementet .
Du är så trevlig .
Åh , Herregud !
Jag pratar inte tyska .
Jag kan inte prata tyska .
Tyskan är inte ett lätt språk .
Pratar du japanska ?
Det här är en japansk docka .
Min hund är vit .
Glöm inte biljetten .
Minns du det ?
Vad är det som saknas ?
Jag brukar diska .
Solen är röd .
På de höstkalla trappstegen upp mot Drottninggatan ligger fimpar bland spridda spottloskor , tillplattade läskburkar och skrynkliga påsar med rester av hamburgare .
I mitt hjärta bor saknaden och längtan efter en annan värld .
Jag har inte sett de någonstans .
Och faktiskt , det var enkelt !
Hon är bara 26 år och driver redan flera bolag .
Hon är en person som kan konsten att vända motgång till framgång .
Och så levde han lycklig i alla sina dagar .
Det var en gång en dvärg som bodde i skogen .
Luciakonserten i Lunds stadshall blev populär .
Betydligt mer än väntat .
800 personer kom för att lyssna på tärnor och stjärngossar .
Boken är också en resa genom 1900-talet .
Åren gick , i makligt tempo och utan att han påverkade världsutvecklingen åt något håll .
Han kom att inse att han gått och blivit gammal .
Det värkte i knäna , alltså levde han nog trots allt .
Att försvara ett fel är att fela igen .
Bara döda fiskar följer strömmen .
En dålig hantverkare klagar på sina verktyg .
Gammal är äldst .
I öknen är sanden billig .
Låt inte vargen vakta fåren .
Man saknar inte kon förrän båset är tomt .
Medan gräset gror , dör kon .
Nöden har ingen lag .
Sovande bonde får drömmande dräng .
Tiden läker alla sår .
Väck inte den björn som sover .
Övning ger färdighet .
Även dåren tros vis om han tiger .
Äras den som äras bör .
Spotta inte i motvind .
Varnad är väpnad .
Varje moln har en silverkant .
Det som göms i snö kommer upp i tö .
Det som göms i snö kommer fram i tö .
Tom är verkligen snål .
En kvinna vars man har dött är en änka .
Vi njöt av att simma i sjön .
Det verkar som att Taro inte har några tjejkompisar .
Tusentals saknas i oväder .
Stormar drabbar sällan området och folk reagerade troligen inte .
Fikonbollarna blir extra snygga om du ringlar lite smält vit choklad över dem när de stelnat !
Jag har ganska stora lår och magrutor , antar att det är muskler , sa hon med ett brett leende .
Vältränade tjejer med god självkänsla är snygga .
Men man får inte banta för mycket .
Älskar du mig ?
Jag heter Hisashi .
Det är en bra idé !
Jag vet att du bor här .
Hon bor i London .
Jag var två gånger i USA .
Jag är student .
Du kan komma med oss om du vill .
En maskerad man i mörka kläder slog sönder två glasmontrar med ett yxliknande föremål .
Flera vittnen som fanns på festen har hörts .
Jag känner mig tom.
Jag behöver köpa en julklapp till min mormor .
De var idel öron när pianisten spelade .
Äppelträden blommar på våren .
Vi har inget socker .
En oskyldig förbipasserande sköts ihjäl mitt på ljusa dagen .
Efter ett gräl med sin fru om bristen på pengar i hushållet rånade en man ett apotek på ett par tusenlappar .
Svenskarna lägger mer på vänsterprasslet .
Ingå i en överenskommelse med mig och bli en ung magisk flicka !
I det mest spännande ögonblicket , såg alla väldigt spända ut .
Åter nås vi av nedslående rapporter om missförhållanden i välfärdsverksamheter .
Det är bara att slå på datorn och nörda loss .
Hon sjunger otroligt bra .
Jag är ledsen , jag tror inte att jag kommer kunna .
Mitt sommarlov är över .
Jag jobbar på McDonalds .
Har inte Jim kommit än ?
Vår skola ligger på andra sidan floden .
Jag är på väg att gå .
Jag trodde att jag skulle kvävas i det överfulla tåget .
Hunden var upptagen med att gräva ner sitt ben i trädgården .
Får jag lämna ett meddelande ?
Har du sett grisen ?
Den tycks ha rymt från stian .
Det var i det huset som jag föddes i .
Det finns ingen slump .
Kvinnan mötte sin mördare av en slump .
När kan jag se dig igen ?
Hon försökte inte att översätta brevet .
Han uppskattar att det nya huset kommer kosta ungefär trettio miljoner yen .
Hon vet bättre än att argumentera med honom .
Min väninna är mycket svartsjuk .
Jag har bara en önskan .
Beyoncé har fött en dotter .
Hans fästmö är redan gift .
Men jag har inga pengar .
Kan du hjälpa mig att översätta dessa meningar till kinesiska ?
Jag kan inte röka .
I allmänhet så är tjejer bättre på att lära sig språk än killar .
Kaniner gillar morötter .
Jag vill dansa .
EU grundas för att få slut på de blodiga krigen mellan grannländerna , som gång på gång hade orsakat så mycket mänskligt lidande och till slut ledde till andra världskriget .
Från och med 1950 börjar en rad europeiska länder samarbeta ekonomiskt och politiskt för att bevara freden .
1950-talet karakteriseras av ett kalla krig mellan östblocket och västmakterna .
Snälla låt mig få plocka upp din syster på stationen .
Jag sprang till min mamma .
Jag lärde mig att cykla när jag var sex år gammal .
Jag kan knappt se utan mina glasögon .
Han drunknade i floden .
Han är den äldsta sonen
Det där rummet är inte stort .
Jag ämnade ringa henne , men jag glömde att göra det .
Jag kom tidigare än vanligt .
Oberoende av vilket instrument du vill lära dig spela , är det viktigaste att inte göra något fel redan i början , ty fel inpräglar sig alltid lättare i ditt minne , än allt som du gör rätt .
Han drack en öl .
Han drack öl .
Vi måste respektera lokala seder .
Koka riset !
De samiska språken hör till ursprungsspråken i Europa och är nära besläktade med de östersjöfinska språken .
Det där verkar vara mycket intressant .
Din dotter är inte längre ett barn .
Skall du presentera mig för henne ?
Jag vill sända detta paket till Canada .
Tom vet inte hur mycket Mary väger .
Picasso målade denna tavla år 1950 .
Kommer hon att kunna lämna sjukhuset nästa vecka ?
Min bror bor i Tokyo .
Yoshio sade att han kan betala upp till 15 000 jen för ett par nya korgbollsskor , men jag anser att det är för mycket .
Vi har en katt .
Vi alla älskar katter .
Det är lättare sagt än gjort .
Jag vill samma svärdet som det !
Igår var han väldigt sjuk men idag mår han mycket bättre .
Vilken sport tycker du mest om ?
Vill du ha påtår ?
Hon log åt mig medan hon sjöng en sång .
Hur firade du din födelsedag ?
Jag vill visa dig hallonbuskarna , lägga ett bär på dina mjuka läppar och öppna dem med en öm kyss .
Fröken Sato är presidentens nya sekreterare .
Jag förstår inte vad du ( vi ) säger .
Allt var väldigt bra .
Jag gav tillbaka kniven som jag hade lånat .
Den där röda tröjan ser bra ut på dig .
Så fort som tjejen såg sin mamma så började hon att böla .
Det gjorde mig ytterst glad .
Hon gillar att prata framför oss .
Jag minns att jag mötte drottningen .
Var snäll och sätt på dig skorna .
Jag antar att du skulle kunna ha rätt .
Varför bestämde du dig för att prata om det nu ?
Ken delade rummet med sin storebror .
Vi har varit gifta i fem år .
Jag sa att jag var förvirrad .
På grund av snön så missade jag tåget .
Jag tror inte att hon skulle förstå det .
Posta det här brevet .
Det är intressant .
Jag behöver inte gå till doktorn längre .
Jag mår mycket bättre .
Jag går hem .
Jag vill dricka en kopp te .
Jag vill inte prata om henne .
Han visste inte vad han skulle göra med den överblivna maten .
Att mingla med folk på fester kan vara förskräckande för blyga människor .
Vad vill du dricka ?
Jag led ett haveri .
Vad betyder katakres ?
Jag steg upp tidigt igår .
Jag mår bra , tack .
Varifrån kommer du ?
Jag är gravid .
Hej då .
Jag behöver en tolk .
Universum hade sin början en torsdag eftermiddag , 13,7 miljarder år sedan .
Var köpte du denne klänning ?
Bomben exploderade för två dagar sedan .
Jag har att skynda !
Han är sjuk .
Han är en hjälte .
Filmen inspirerades av boken med samma titel .
Många har samlats .
Tom ville inte göra något han skulle komma att ångra .
Mary gillar att festa .
Det verkar som att Mary är full igen .
Måste jag hålla ett tal ?
Mary försökte trösta Tom .
Jag sov som en stock .
Mary kände sig utstött .
Depression är vanligt bland unga vuxna som har Asperger syndrom .
Jag beställde nya möbler .
Vad pratar hon om ?
Regniga dagar gör mig deppig .
Finns det en bank i närheten ?
Han har blivit längre och längre .
Jag såg filmen fem gånger .
En änka är en kvinna , deras make har dött .
Vem äter bin ?
En otrevlig känsla är aldrig bra .
Sanningen kommer fram när förstånd och känsla stämmer överens .
Han emigrerade till Australien .
Koranen som jag har är tvåspråkig , den är tryckt på arabiska och esperanto .
Tillsvidare har jag varit i mer än tio främmande länder .
Kommer du att delta i festen ?
Runt staden rinner en flod .
Runt staden flyter en flod .
Landet förklarade krig mot sitt grannland .
Jag har inte sett henne på länge .
Jag skojar inte .
Hur länge tar det till fots ?
Vill du att jag skall koka kaffet ?
Polisen talade med en man på gatan .
Tjänarinnan höll redan på att städa rummet när Carol kom in .
Han stack handen i fickan och letade efter sin plånbok .
I begynnelsen var ordet .
Var det ett nyord ?
Hon strykte sin skjorta .
Hon gav oss ett inexakt svar .
Han blev en mycket god musiker .
Så länge man har ett mål , finns det hopp .
Utsvultna och vanskötta duvor omhändertogs .
Duvorna var innestängda utan mat i ett smutsigt utrymme.Två hade hunnit dö .
Jag skämtar inte .
Jag spelar Sudoku då istället för att fortsätta störa dig .
Han är på sjukhuset .
Tom är en främling i den här staden .
Nuförtiden verkar alla vara lyckliga .
Du borde ha bett om ursäkt till henne .
De skrattade åt min idé .
Jag skulle vilja simma i den här floden .
Det är möjligt att Jane inte är hemma just nu .
De började sälja en ny typ av bil i Tokyo .
Jag har spenderat mycket pengar på mitt hus .
Jag ser fram emot att träffa dig .
Tom vet inte vart han skall gå .
En sjukdom förhindrade honom från att gå ut .
Fram tills förra veckan hade jag inte fått något svar .
Det var inga varningar överhuvudtaget .
Den korta kvinnan har på sig en svart kostym .
Allt i denna värld är blott en dröm .
Problemet är att vi inte har någonstans att vara ikväll .
Ett hundra cent blir en dollar .
Du är längre än mig .
Jag kommer inte ihåg ditt namn .
Gå upp tidigt på morgonen .
Den här bussen får plats med femtio personer .
Vi tittade alla ut genom fönstret .
Jag antar att han kommer tillbaka snart .
Vad är det för skillnad mellan en by och en stad ?
Gillar du att äta fisk ?
Han kommer kunna gå upp och gå om ungefär en vecka .
Han berättade sin livshistoria för mig .
Han tjänar tre gånger så mycket som jag .
Han la boken på hyllan .
Du borde inte säga såna saker när barn är i närheten .
Du ser precis ut som din storebror .
Du går inte upp lika tidigt som din syster , eller hur ?
Vart i Turkiet bor du ?
Hon hade precis börjat läsa boken när någon knackade på dörren .
Vilka språk talas i Amerika ?
Det där är anledningen varför han blev arg .
Det där är varför han blev arg .
Kaniner har långa öron och korta svansar .
Om inte den där gitarren vore så dyr , så skulle jag kunna köpa den .
Jag sa till henne en gång för alla att jag inte skulle gå och handla med henne .
Jag är överraskad att du vann priset .
Hon kommer förmodligen .
Det är ungefär lika stort som ett ägg .
Det är väldigt varmt idag .
Klockan är redan elva .
Jag skjuter upp min resa till Skottland tills det blir varmare .
Jag vet inte exakt när jag kommer att komma tillbaka .
Jag kommer tillbaka snart .
Hon är nyfiken på att få reda på vem det var som skickade blommorna .
Hon vill veta vem det var som skickade blommorna .
Håll bollen med båda händerna .
Jag är på åttonde våningen .
När man har fått in en dålig vana , så är det inte enkelt att bli av med den .
Jag kan inte komma ihåg den låtens melodi .
Han visade mig en massa vackra bilder .
Hon hjälpte den gamla mannen över vägen .
Jag behöver gå ner i vikt , så jag håller på med en diet .
Vargar brukar inte attackera människor .
Han återvände hem efter att ha varit borta under tio månader .
Vill ni att jag skall koka kaffet ?
Vill ni att jag skall koka kaffe ?
Kärleken är blind .
Kontakta henne om du har några frågor .
Vi har gått runt hela sjön .
Hon har inte varit i skolan på fem dagar .
Det är svårt att förstå hans teori .
Det är upp till dig att bestämma om vi skall gå eller inte .
Han är tre år äldre än henne .
Hon håller på med en diet .
Det verkar som att jag har en lätt förkylning .
Rätta mig om jag har fel .
Jag är nyfiken .
Jag är rädd för hundar .
Jag har en massa arbete att göra imorgon .
Han är DJ .
Jag har levt här under en lång tid .
Jag har en känsla av att hon kommer att komma idag .
Det kommer inte att fungera .
Hon skadades i en bilolycka .
Hur kommer det sig att du alltid är sen ?
Jag tycker att det är tragiskt att inte ha några vänner .
Jag översatte dikten så gott som jag kunde .
Jag kände mig väldigt lättad när jag hörde nyheterna .
Jag är säker på att jag kommer vinna tennismatchen .
Jag höll i repet hårt så att jag inte skulle falla .
Jag kunde inte gå på hans födelsedagskalas .
Jag kommer aldrig att glömma din vänlighet .
Jag uppskattar verkligen din vänlighet .
Jag tyckte att den här filmen var väldigt intressant .
Jag dricker alltid två koppar kaffe varje morgon .
När jag kom hem , upptäckte jag att jag hade tappat bort min plånbok .
Oavsätt hur mycket hon äter , så går hon aldrig upp i vikt .
Det han sa visade sig vara en lögn .
Hur länge kommer det här kalla vädret att hålla på ?
Hur länge kommer det här kalla vädret att fortsätta ?
Jag kommer känna mig ensam när du har gått .
Hur lärde du dig att spela fiol ?
Han är vänligt mot alla sina klasskamrater .
Han kunde inte komma tillbaka , då han var sjuk .
Han var sjuk , så han kunde inte komma .
Hans försök med att simma över floden misslyckades .
Han lät mig sova över en natt .
Han gillar verkligen musik mycket .
Han älskar musik .
Han gillar musik mycket .
Han kan inte ha sagt något så dumt .
Prata inte runt den heta gröten , säg det genom blommorna .
Han tappade greppet om repet och föll ner i floden .
Jag tycker att hon är en ärlig kvinna .
Jag kommer att vara sexton år gammal på min nästa födelsedag .
Låt mig berätta för dig om fallet .
Jag kommer förklara incidenten .
Jag ville ringa några telefonsamtal .
Jag har hört den franska versionen av den här låten .
Jag har hört den låten sjungen på franska .
Jag är inte säker på när han kommer att komma .
Jag tror att jag skall köpa en ny bil .
Premiärministern kommer att hålla en presskonferens imorgon .
Hur hände trafikolyckan ?
Han har vanan att läsa tidningar under måltider .
Han övar på att spela gitarr tills sent på kvällen .
Han gick vilse när han var ute och gick i skogen .
Han försökte att göra sin fru lycklig , men han kunde inte .
Han gick ut ur rummet utan att säga ett ord .
Han gick in på banken utklädd som en vakt .
Han älskar att resa .
Han gick ut ur rummet så fort som jag gick in .
Det finns ingen chans att han kommer att återhämta sig .
Han har ingen chans att återhämta sig .
Han sover under dagarna och jobbar under nätterna .
Han visade mig hennes fotografi i smyg .
Han visade mig hennes foto i smyg .
Han visade mig hennes bild i smyg .
Han verkade besviken över resultaten .
Han litar mycket på sin assistent .
Han studerade hårt så han inte skulle misslyckas .
Han har ett stort hus och två bilar .
Han gick långsamt så att barnen skulle kunna klara av att följa efter .
Han gick långsamt så att barnet kunde följa med .
Vi skulle vilja beställa 18 ton olivolja .
Av misstag svängde han vänster istället för höger .
Vi åker och fiskar då och då .
Faktum var att han till och med älskade henne .
Flygplan kan höras långt före de syns .
Ett spädbarn sover i vaggan .
Var snäll och stäng dörren efter dig .
Tom ser Mary som en hjältinna .
Förlåt , det var inte min mening att sparka dig .
Det här är det värsta av allt .
Hallå där !
Din baseboll hade just sönder mitt fönster .
Vi kan inte vara utan vatten ens för en dag .
Min cykel behöver lagas .
Har du skrivit upp telefonnumret ?
Har du skrivit ned telefonnumret ?
Hon ger sin son för mycket pengar .
Hon läser tidningen varje morgon .
Han talade inte såvida han inte blivit tilltalad .
Läraren underströk vikten av att föra anteckningar .
Kan du sänka priset till tio dollar ?
Jag vet inte hur man spelar golf överhuvudtaget .
Jag tycker att han är skicklig .
Jag tycker att han är en skicklig person .
Jag var inte medveten om att du mådde så dåligt .
Jag tycker att du borde tänka på framtiden .
Jag tycker att du behöver tänka på framtiden .
Jag gjorde ett allvarligt misstag på provet .
Jag gjorde ett dåligt misstag på provet .
Jag lånade ut en del pengar till min vän .
Ofta kommer han inte till skolan .
Det var inte nödvändigt att han skulle ta med ett paraply .
Han behövde inte ta med sig ett paraply .
Han tänkte att det skulle vara vettigt att acceptera erbjudandet .
Han är väldigt smart , så alla gillar honom .
Han säger alltid elaka saker om sin fru .
Bäckens porlande musik smeker apelsinträdens blad .
Cowboy hoppade snabbt ut genom fönstret .
Idag , den 6 februari , är det den samiska kulturens dag , samernas nationaldag .
Är han en lärare ?
Hon är envis .
I Sameland talar man många språk .
Minns du den än , minns du den lyckliga tiden ?
Är mjölken god ?
Mannen bad mig om litet pengar .
Han betraktade himlen .
Tatoeba har inte alla språk som jag behöver .
De är en finländsk , svenskspråkig grupp .
Vi behöver fler arbetare .
Arbetarna var stolta över sitt arbete .
Jag är älskad .
Jag kommer att bli älskad .
Jag var älskad .
Jag skulle vara älskad .
Var älskad !
Hon befann sig på platsen för brottet .
Hon var på brottsplatsen .
Du skall bli tvättad .
Ni kommer att bli tvättad .
Man kan inte ha framgång om man inte arbetar mycket .
Man kan inte vara framgångsrik ifall man inte jobbar mycket .
Varför är himlen blå ?
Vad vet du om näringslivet i Sverige ?
Det är ingen leksak !
Min mor är arg .
Pojken köper en hund .
Jag känner mig gammal .
Jag är van vid att äta ensam .
Jag fick ett erbjudande jag inte kunde motstå .
Han har en utländsk bil .
Jag än inte alls intresserad av politik .
Jag har en god idé .
Var inte ett sådant arsle !
Katten har sovit på bordet .
Vem är det som spelar gitarr ?
Jag har två döttrar .
En fånge rymde från fängelset .
Vi såg en skymt av slottet från vårt fönster i tåget .
Vita duvor är vackra fåglar .
Vi bor inte i länder , vi bor i våra språk .
Det är ditt hem , där och ingen annanstans .
Varför trodde du inte på mig ?
Vem är det som sover i min säng ?
Jag har bestämt mig för att berätta för honom att jag älskar henne .
Pilen missade sitt mål .
Vad påminner denna hatten dig om ?
Latin är ett dött språk .
Det är ett foto av en apa i samband med apans år .
Han gav inte ett enda ord till svar .
Enligt tidningen var det ett jordskalv i Peru .
Det var 1912 som Titanic sjönk under sin första resa .
Han är strax över trettio .
Hon hittade ringen som hon hade tappat under resan .
Han är hennes vän .
Guldpriset ändras dagligen .
Jeans är mode bland flickor nu för tiden .
Han liknar sin far .
Han liknar sin pappa .
För att säga det rakt ut ; Jag gillar inte honom .
Läraren har rätt .
Jag råder dig att åka hem .
Jag besöker dig nästa söndag .
Jag ser på tv varje dag .
Jag har tappat min börs .
Hon äter inte kött , eller hur ?
Det är ett simpelt fel .
Först i går fick vi reda på det .
Jag är en människa med många fel , men det är fel som enkelt kan rättas till .
Vi uppskattade skadan till tusen dollar .
Jag öppnade asken .
Den var tom.
Vem är din kinesiskalärare ?
Det är dags att gå och lägga sig .
Vilken del av Kanada kommer du ifrån ?
Hon gifte sig vid en ålder av sjutton .
Jag är mycket intresserad av fotboll .
Vi har talat om er .
Problemet är att jag inte har några pengar på mig .
Columbus upptäckte Amerika 1492 .
Vad gör du för att få tiden att gå ?
Han ändrade plötsligt sin inställning .
Böterna ska betalas kontant .
Jag har bott i Koenji .
Mitt rum är mycket litet .
Jag försöker gå ner i vikt .
Kom hit !
Kylie Minouge är den bästa sångerskan jag någonsin har sett !
Han bor utanför stan .
Min katt dödade denna musen .
Det påstås att det snart kommer ett val .
Planen stöddes av praktiskt taget alla närvarande .
Skolan är på gångavstånd från mitt hus .
Tom gick vilse .
Vi är lika inför lagen .
Vilken är din favoritprotestsång ?
Hon beordrade honom att städa upp sitt rum .
Han längtar efter stadsliv .
Flickan var snäll och berättade vägen till museet .
Det är ingen tvekan om vem som blir vald .
Det står bra till med min familj , tack .
Min familj mår bra , tack .
Han erkände att han hade tagit mutor .
Japan behövde kontakt med västerlandet .
Min bror kan komma att behöva en operation för knäskadan .
Hunden följde mig .
Jag är glad att se dig !
Hon brukade gå upp tidigt .
USA är en republik medan Storbritannien inte är det .
Hon är inte doktor .
Jag är inte rädd .
Rie och jag har gått i samma skola .
Jag tycker du har blivit mycket bättre på engelska .
Du kan välja antingen det ena eller det andra .
Jag går upp i vikt , för jag äter mycket godis .
Var är den vackraste platsen i världen ?
Tom är lika lång som Jim .
Önskar ni att ni var rika ?
Det är vackert väder idag .
Har du en speciell meny för vegetarianer ?
De här blommorna är vackra , inte sant ?
Får man fotografera i detta huset ?
Det är inte alla fåglar som kan sjunga .
Jag är stolt över dig .
Oavsett hur mycket jag försöker kan jag inte komma på hennes adress .
Oavsett hur mycket jag försöker kan jag inte komma ihåg hennes adress .
Jag har två bröder och en syster .
Vanligtvis äter vi tre gånger om dagen .
Du förväntar dig för mycket av henne .
Varför kom du inte ?
Försök att se det som det är .
Försök att se saken som den är .
Tack för informationen .
Jag har en vän vars far är lärare .
Jag har en vän vars pappa är lärare .
Nancy vill ha ett par röda skor .
Ledarhundar hjälper personer som inte kan se .
Har ni julledigt i Japan ?
Den nya tunneln kommer att förbinda Storbritannien med Frankrike .
Island hörde till Danmark .
Fåglar sjunger tidigt om morgonen .
När inträffade händelsen ?
Var snäll och sitt kvar .
Jag tyckte det var en bra bok , men Jim hade en annan uppfattning .
Trädgården var full av vackra blommor .
Den här klänningen kan se lustig ut , men jag gillar den .
Det är några båtar i sjön .
Biblioteket ligger mitt i stan .
Om du älskar mig , älska också min hund .
Hon brukade dricka öl .
Vi ogillar regnet .
Förra månaden gifte hon sig med Tom .
Filmen började klockan 2 .
Han köpte ett par nya handskar .
Se på huset med det röda taket .
Han ser inte ut som en intelligent pojke .
Hon går på en diet .
Jag vill veta detaljer .
Den mannen dog av lungcancer för en vecka sedan .
Den kvinnan har två väskor .
Taro , vill du vara så snäll och hjälpa mig ?
Han knackade på dörren .
I går var det fredag och i övermorgon är det måndag .
När jag blir stor ska jag bli kung !
Det är ofarligt att äta fisken .
Han bor sex hus från mig .
Inget saknas .
Mm-hm .
Det tror jag med .
Han gillar att se på tv .
Jag är inte din docka .
USA är en republik .
Vi gifte oss för sju år sedan .
Den boken säljer bra .
Kom du med tåget ?
Rom byggdes inte på en dag .
Han la handen på min axel .
De böckerna tillhör min syster .
Folk är rädda för krig .
Ingen visste det .
De har ännu inte fastlagt datumet för sitt bröllop .
Jag vet inte exakt när jag kommer tillbaka .
De tolv stjärntecknen är : Väduren , Oxen , Tvillingarna , Kräftan , Lejonet , Jungfrun , Vågen , Skorpionen , Skytten , Stenbocken , Vattumannen och Fiskarna .
Var såg du de här kvinnorna ?
Gör dig inget besvär !
Hur har din fru det ?
Vädret blev bättre .
Mjölk håller inte länge när vädret är varmt .
Var var du på din semester ?
Var snäll och ge mig ett glas mjölk .
Vad sägs om att spela tennis på lördag ?
jag ser fram emot att se dig till jul .
Är katten på stolen eller under den ?
Vill du ha något att dricka ?
Min vän gjorde slut med sin flickvän och nu vill han gå ut med mig .
Jag fann honom extremt intelligent .
Det retar mig att de har glömt att betala .
De äpplena är stora .
Jag går ut och leker .
Följer du med ?
Du borde ha hållit det hemligt .
Vin hjälper matsmältningen .
Efter oss syndafloden .
Jag hårdkokte ett ägg .
Jag började studera esperanto när jag var i tonåren .
Kan du springa fort ?
Hon har få vänner .
Jag har hört nyheten om att det har varit en stor jordbävning i Awaji .
Räkna från ett till tio .
Män är svin .
Han dog i cancer förra året .
Hon röker 20 cigaretter om dagen .
Han uppför sig som ett barn .
John har en bil från Japan .
Gick du upp sent ?
Jag gav tiggaren alla pengar jag hade .
Jag kommer att vara där i morgon .
Du måste läsa mellan raderna .
Han tog ledigt en vecka .
Är han fortfarande kvar ?
Min mor går på diet .
Min mamma går på diet .
En ny filial öppnar i Chicago nästa månad .
Han har blont hår .
" A " är alfabetets första bokstav .
Jag vill gärna träffa Er igen i nästa vecka .
Du kan inte ha förstått vad han sa .
Det är gratis .
Jag tror att den här medicinen kan hjälpa mot din sjukdom .
Går din klocka rätt ?
Hur har du det ?
Den dunkudden ser dyr ut .
Man har ljugit för dig .
Han måste älska dig .
Vem ritade det ?
Vad står det skrivet på trafikmärket ? -Enkelriktat .
Jag är tvungen att hitta ett deltidsarbete .
Mor köpte en vacker kjol till mig i söndags .
Jag tänkte på dig .
En dator är en komplex maskin .
Jag är väldigt glad över att träffa dig .
Det var en jordbävning i går .
Kom inte för nära mig .
Jag är förkyld .
Jordbävning kan inträffa när som helst .
De blommorna växer i varma länder .
Vi kommer att vänta på dig där .
I dag är det årets varmaste dag .
Hon log .
I morgon är det jul .
Du gör mig besviken .
Jag står till ditt förfogande .
Är de här nyheterna sanna ?
Korta brev och långa vänskaper , det är min devis .
På marken lever olika insektsarter .
Ursäkta , hur sent är det ?
Där är en katt i köket .
Det är bara två veckor till jul .
Varje stad i USA har ett bibliotek .
Jag läste brevet för honom .
Vi har precis fått information om att fienden ligger i bakhåll på vägen två mil längre fram .
Soldaten slog samman klackarna .
Efter vintern kommer våren .
Det som ser enkelt ut vid första ögonkastet visar sig vara svårt .
Hur mycket har du betalt för dem ?
Ibland går jag till arbetet och ibland cyklar jag , eftersom jag bor mycket nära arbetet .
Chips är inte bra för din hälsa .
Nyfikenhet dödade katten .
Byborna bygger en träbro över floden .
Min lärare är herr Haddad .
Hon vill bli simultantolk .
Tåget har inte kommit ännu .
Gör som läkaren sagt .
Har du någonsin varit i utlandet ?
Det var tur i oturen att ingen dog .
Åh !
Min dator är trasig .
Herr Kinoshita glömde sina glasögon på kontoret i går kväll .
Han tog på sig den svarta överrocken .
Jordens måne är en naturlig satellit .
Tom har tre onklar .
Om du vill hitta den sanna vägen , måste du liksom sköldpaddan hitta balansen mellan det som är hårt och det som är mjukt .
Jag läste att Brasiliens president är en kvinna .
Hon kallas Dilma .
Bara för att du inte finns på riktigt så betyder det inte att du kan säga åt mig vad jag borde göra .
Berätta en zombie historia för mig .
Burj Khalifa är världens nuvarande högsta skyskrapa .
Jag behöver köpa frimärken .
Jag kommer aldrig att lämna dig .
Moder Teresa föddes 1910 i Jugoslavien .
Var är ingången ?
Jag talar inte kinesiska .
Elbrus är Europas högsta berg .
Jag betalar med mitt kort .
Han dömde Brown till hängning .
Jag har slutat med öl .
Var snäll och stäng av motorn .
Vi förknippar namnet Darwin med evolutionsteorin .
Jag måste vara hemma vid tio .
Jag kan inte höra dig , vänligen tala högre .
Har du böcker på esperanto ?
Jag vill kunna läsa japanska .
Det finns inga matbutiker i närheten .
De sårade kom med ambulans .
Staden var öde .
Livet är orättvist .
Hans skjorta var grå och slipsen gul .
Han har god anledning att tro det .
Jag tar den gula .
Men det var förstås länge sedan .
Han kände i fickan efter tändaren .
Den här ölen har hög alkoholhalt .
Han hade i arbetet kommit i kontakt med några utlänningar .
Min vän George ska till Japan i sommar .
Jag behöver nycklarna .
Lägg inte dina grejer i gången .
Låna aldrig en bil .
Jag kände mig lätt som en fjäder .
Vi träffades en vinter .
Räcker tiotusen yen ?
Jag börjar så sakta tycka om Ken .
Han har inte lyckats än .
Hon ser ung ut för sin ålder .
Du borde äta mer frukt .
Här kommer vår lärare .
En 90-gradig vinkel kallas en rät vinkel .
Harry är bara 40 .
Välkommen hem till oss !
Välkomna hem till oss !
Vilken är din favoritsvordom ?
Det finns ett akut behov av bloddonationer .
En ung flicka satt vid ratten .
Dagen gryr .
Jag måste ta ett paraply med mig .
Du borde komma och hälsa på oss !
Ni borde komma och hälsa på oss !
Och så förälskade sig lejonet i tackan .
Alla pratade om det .
Dubbelklicka på ikonen .
Jag frågade honom vad han hette .
Håller isen ?
Jag läser den här boken .
Den här kniven är för slö för att skära med .
Boten skall betalas i kontanter .
Jag hatar när mina kläder luktar cigarettrök .
Det här ägget är färskt .
Medtävlanden tjuvstartade två gånger .
Får jag titta på tv nu ?
Krig är fred .
Frihet är slaveri .
Okunnighet är styrka
Du är guld värd .
Vi träffas här en gång i månaden .
Vatten består av syre och väte .
Jag kunde hjälpa henne .
Idag är det imorgon vi oroliga igår .
Japans huvudgröda är ris .
Vi måste ta itu med det här problemet .
Jag fattar .
Hon kom inte innan två .
Titta inte ut genom fönstret .
Vems rum är det här ?
Jag lärde känna honom när jag var student .
De hämtar våra sopor varje måndag .
Mayuko verkar klok .
Hur skiljer sig din åsikt från hans ?
Hon blir sen till maten .
Jag avskyr att ha med kräsna barn att göra .
Jag var på väg ut .
Behöver du hjälp med att bära något ?
Pojken gick vilse i skogen .
Oavsett hur snabbt du kör hinner du inte dit i tid .
Han berättade inte för John om olyckan .
Han hjälper inte till hemma .
Vi skulle samarbeta i projektet .
Jag sitter och studerar på biblioteket .
Jag går och tar ett glas öl .
Du känner , det är sant .
Jag väcker på morgonen vid halv sju .
Teatern är tråkig .
Vill du komma att gå och shoppa ?
Där kan man äta mycket bra .
Nästa artisten är fantastisk .
Hans mobil har blivit stolen .
Jag vilja flytta på Australien .
Vill du sova hemma hoss mig ?
Det är din först arbetsuppgift .
Tom måste erkänna sitt lagbrott .
Jag vill inte gå ut .
Är det vad du vill ?
Jag älskar filmar .
Han är på tåget .
Alice har fantastiska benen .
De kom inför er .
Blunda och sov .
Hur länge har de varit här ?
Jag tror inte det blir bättre än så !
Kejsar Hadrianus lät bygga Hadrianus mur .
Han förlorade hans nya klocka .
Rör det inte !
Jag gick an om .
Matchen slutade utan malen .
Jag har satt på TV och man uppträdde Grand Prix .
Mannen vaknar .
Hon har en viktig roll i vår organisation .
Mina skor måste lagas .
Varför kommer hon inte ?
Nu är jag ryckigt trött .
Jag behöver en cigarett .
Ska vi fika ?
Det är inte en bra idé .
Jag tar en promenad .
Jag skulle vilja förbättra min franska , men Jag får inte tid med .
Har du tid att äta middag med mig ikväll ?
Det är inget att bry dig om .
Vattenverket ligger inte långt från mitt hem .
Jag är dålig på tennis .
Jag fick syn på pojken .
Jag hann dit i tid .
Jag måste ha drömt det .
Jag har varit hos tandläkaren .
Tom visste inte var han skulle börja .
Han tycker om att simma .
Vad är det för fel på mig ?
Han förklarade sin situation för mig .
Kan du släcka ljusen ?
Kan du släcka stearinljusen ?
Han valdes till president .
Jag skiter i vad du säger !
Tom var klädd helt i svart .
Tom räddade hunden ifrån att bli uppäten av de hungriga soldaterna .
Jag skakade hand med Jane .
Vad är haken ?
Det erbjudandet låter för bra för att vara sant .
Vad är haken ?
Några av mina klasskamrater gillar volleyboll , medan andra gillar tennis .
Det är en genant sjukdom .
Jag svettas varje dag .
De analyserar proven .
Hon försvann utan papper .
Blond tjejen har mycket bra bröst .
Vem dödade henne ?
Svaret är inte korrekt .
Det finns inget mer salva .
Söndags matchen ska bli avgörande .
Ingenting är lätt .
Du är tokig !
Bilal gick i skolan .
Mina läppar är stängt .
Jag har sett Liz i morse .
Hon är gammal .
Det zoo äger två okapi .
Jag har hört ingenting .
Vi är man och fru .
Vägarna är lortig .
Här kan ni röka .
Det är hans julklapp .
Han satt alldeles tyst och tittade rakt fram .
De körde igenom flera samhällen på vägen .
Hon tittade på alla hus som gled förbi .
Hon undrar hur det se ut där de skulle bo .
Men allra mest undrade hon vad hette henne .
Då är jag framme .
Nå vad tycker di om mig ?
Han lastade ur bilen .
Hon stängde försiktigt ytterdörren .
Så bullrig det var därinne .
Rummet verkar väldigt mörkt och kusligt .
Hon kände sig plötsligt så liten .
Det ekade ödsligt .
De gick uppför trappan .
Jag letade efter mitt rum .
Du ska hitta dina leksaker och böcker .
Jag kände mig genast lite bättre .
Vad är det för filtillägg ?
Hon kan spela den här melodin på piano .
Nyheten om hennes död kom som en blixt från klar himmel .
Vad gör tvättbjörnen i köket ?
Liljorna som täcker den blå dammen hindrar mig från att se min avbild i vattnet .
Transformation är födelse och död på en och samma gång .
Glöm aldrig den skatt som finns i djupet av din själ : medkänslans milda flamma som gör varje dag meningsfull .
Ingen förstår mig .
Jag talar inte japanska .
Vi har en kvadratisk tabell .
Tystnad är guld .
Frankrike är i Västeuropa .
Envar har rätt till skydd för de moraliska och materiella intressen , som härröra från varje vetenskapligt , litterärt eller konstnärligt verk , till vilket han är upphovsman .
När registrerade de medlemmarnas namn ?
Geologen klev in i limon .
Jag köpte inte den där boken .
Du är i bättre form än jag .
Kristus är uppstånden !
Han är min vän .
Var ligger Mississippi ?
Tom är inte här .
Mari och Maki är systrar .
Alla vill träffa dig .
Du är känd !
Han är alltid väldigt artig .
Varför går inte människor i ide ?
Du har två bollar .
Du har två kulor .
Det här gräset behöver klippas .
Vi måste försöka bryta dödläget .
Snart är det din tur , Bashar !
Har du hört av henne ?
Kenya blev självständigt 1963 .
När han kom hem , sov barnen redan .
Vem sjunger den här sången ?
De här grejerna är inte mina .
De här sakerna tillhör inte mig .
Får jag göra nånting ?
Han satt där för att röka en pipa .
Varför tittar du på mig på det där sättet ?
Han tycker inte om fisk .
Jag tror på vad han säger .
Har du redan tagit din medicin ?
Jag tror på honom .
Hur lat är du egentligen ?
Han snarkade högt medan han sov .
Du ska dit utan meg .
Min syster är mycket klok .
Min faster har tre barn .
Min moster har tre barn .
Jag vill titta på filmen .
Får jag komma med ?
Får jag vara med ?
Jag har svarta ögon .
Jag träffade en hund på vägen hem .
Min mor är alltid upptagen .
Jag skulle vilja gärna betala .
Jag är trött på läxor .
Du behöver inte säga upp jobbet .
Jag älskade att läsa då jag var liten .
Jag är mycket trött .
I vilken klass går din lilla syster då ?
Det kan jag inte tro på .
Vi ska segla till Danmark .
Det är svårare än vad du tror .
Det här äpplet smakar dåligt .
Ge mig mina glasögon .
Jag har sovit , och du ?
Ett år har tolv månader .
Ska vi till bio ?
Jag tycker om regn och snö .
Han är en modern pojke .
Jag mår bra .
Läraren och eleverna är i museet .
Tvätta dina fötter .
Jag är ingen läkare .
Mina barn är i skolan .
Det var en gång en kung som hade tre döttrar .
Jag ska bygga en stor byggnad .
Jag behöver hjälp .
Jag ska skriva en bok .
Jag är gammal .
Ingen översätter mina satser .
Jag är glad .
Hur mycket pengar har du ?
Hur många pengar har du ?
Jag måste se det !
Många människor pratar bara ett språk .
Jag hoppas inte .
Katten har två öron .
Jag skulle vilja växla pengar .
Jag har ingen bil .
Jag vill gifta mig med honom .
Jag sjunger nu .
Katten har nästan blivit påkörd av en lastbil .
Den här engelska boken är för svårt för mig att läsa .
De här böckerna tillhör dem .
Dessa böcker är deras .
Han lyssnar på allt vad du säger .
Hela världen tittar på oss .
Vår skola är åttio år gammal .
Allt lyses av solen .
Han kommer tillbaka klockan fyra .
Tyvärr Nancy hade rätt .
Hennes enda fritidsintresse är att samla på frimärken .
Han är sitt vanliga jag .
Skala äpplet innan du äter det .
Vad är populärt nu ?
Vad är inne nu ?
Vad är på modet nu ?
Är du rädd för skräckfilmer ?
Är du rädd för rysare ?
Det är lättare att lyfta än att landa .
Jag vill dricka något kallt .
Paris är en ganska dyr stad .
Tom har bevisat att det fungerar .
Tom har bevisat att den fungerar .
Tom har bevisat att det går .
Varför var du där ?
Min bil är stor nog för fem personer .
Han har nått sitt mål .
Min familj är inte så stor .
Skolan börjar den åttonde april .
Han var upptagen .
Jag älskar att promenera ensam .
Tom tittar för mycket på tv .
De bestämde sig för att bygga en bro .
Stjärnorna blinkade på himlen .
För mig är det viktigt .
Jag bodde i Tokyo för nägot är sedan , men nu bor jag i Kyoto .
I går var jag för sjuk för att gå till skolan .
Vi är inte i fara nu .
" Mina tänder är för svaga för att äta ett äpple " sa pojken .
Vet du vad det betyder ?
Jag har ont i tanden .
Ja , jag tycker om det .
Han hugger träd uppe på fjället .
Var så god och ge mig något att äta .
Min dröm är att studera utomlands .
En kungs dotter är en prinsessa .
Jag somnade framför TV-en .
Jag har ätit gott .
Gissa vem som kommer i kväll .
Jag skulle hellre vara en fågel än en fisk .
Får jag äta ?
Jag har byggt ett nytt hus .
Tack för senast .
Mina föräldrar älskar varandra .
Hon ringde sin mor .
Hon kom hem sent på kvällen .
Jag har inte någon bil .
Vems vän är du ?
Jag har skrivit ett brev .
Han är min lärare .
Får jag gå nu ?
Den här bron byggdes för två är sedan .
Vad säger han ?
Ni måste hem .
Du måste hem .
Vi har inte sett nånting .
Hon spelar piano varje dag .
Min mor är inte hemma .
Min mor är ute .
Jag kan spela gitarr .
Weigongcuns tunnelbanestation har tre utgångar .
Ett kuvert och ett frimärke , tack .
Flickan gick till skogen för att plocka svamp .
Du får komma med .
Jag vet .
Han bor i Osaka .
Du äter ingenting .
Om du inte äter dör du .
Jag ser ingen .
Bättre en fågel i handen än tio i skogen .
Det här är huset som min farbror bor i .
Han mår bra .
Det är kallt idag .
Vinden blåser från öst .
Han tog henne i handen .
Jag har ingen tid nu .
Krokodilarna har vassa tänder .
Hon säger hon tycker om blommor .
Vad gör din son ?
Den här fågeln kan inte flyga .
Är du tio ?
Är du tio år gammal ?
Jag ringer dig om en timme .
Jag går till parken .
Jag ska till parken .
Den är vit som snö .
Jag vet att du är rik .
Vilken tid kan du komma ?
Maria har långt hår .
Min bror är inte så stor som jag .
En hund har bitit mig i benet .
Han ska följa min råd .
Vem kommer med mig ?
Han drack tre glas vatten .
Jag gick till stationen .
Vi är båda studerande .
Var har du köpt de där skorna ?
Jag tuggade tuggummi .
Jag har inga pengar men jag har drömmar .
När kommer du ?
Jag vill inte att du berättar det för henne .
Du behöver inte svara på de här frågorna .
Jag vill skriva en bok .
Jag ville dit .
Hur länge ännu , Catilina , skall du missbruka vårt tålamod ?
Den unga mannen är läkare .
Jag är höjdrädd .
Gör honom inte besviken .
Ta seden dit man kommer .
Jag är inte alls trött .
Fisken är .
Hämnd är den bästa hämnden .
Om du verkligen vill lyckas måste du tycka om att äta gift .
Om du är rädd för att dö har du redan dött .
Han satt där med sina ögon stängda .
Den tillhör min bror .
Japan är ett vackert land .
Fortsätt träna när du fått lite te i dig .
Du borde koncentrera dig på vägen när du kör .
Drick medicinen .
Våra gudar är döda .
Talar du klingonska ?
Jag kan inte klingonska .
Qo ' noS är klingonernas hemplanet .
Jag talar klingonska med dig .
Fyratusen meningar kan översättas på ett år av en talande man .
Har du inga pengar så får du klara dig utan .
Han dog en ärorik dysenteridöd .
Jag tror inte att det kommer att regna i eftermiddag .
Vi har tre flygplan .
Kjolen är grön .
Jag blöder om knät .
Jag tittade på matchen från början till slut .
Bland hans musikaliska verk finner man tolv operor och operetter .
Ser man på !
Jag behöver kaffe .
Herre , var nådig mot min son , ty han är epileptiker och lider fruktansvärt därav , för han faller ofta in i elden , och ofta ner i vattnet .
Elden är utan nåd .
Elden har ingen nåd för någon .
Kapitulera eller dö !
Köp eller dö !
Hon är gammal nog för att resa själv .
Jag beter mig inte som du .
Gör som jag !
Jag kommer inte ihåg deras namn .
Jag kommer inte på vad de heter .
Han spelade golf varje dag under semestern .
Sin älskades doft känner man alltid .
Fira !
Imorgon ska vi kanske dö !
Jägaren gör inte det liggande bytet sällskap .
Det där var en utmärkt putt .
Esperanto talas i 120 länder runt om i världen .
Visst är det möjligt om man vill .
Du vänjer dig snart vid din nya skola .
Vad betyder " Tatoeba " ?
Ty mörkret har passerat , och legenden gror ännu .
Det betyder slutet för ondskan , och för alla fiender av Skyrim .
Jag säger er , jag säger er , den Drakfödde kommer !
Kossan säger " mu " , tuppen säger " kuckeliku " , grisen säger " nöff , nöff " , ankan säger " kvack , kvack " och katten säger " mjau " .
Kossan muar , tuppen galer , grisen grymtar , ankan kvackar och katten jamar .
Tuppen galer " Kuckeliku ! " om morgonen .
Tuppen pickar på mitt ben .
Var ligger den svenska ambassaden ?
Var finns det en svensk ambassad i USA ?
Det finns en svensk ambassad i Washington D.C.
Var ligger den franska ambassaden ?
Var ligger den tyska ambassaden ?
Var ligger den kinesiska ambassaden ?
Var ligger den australiska ambassaden ?
Var ligger den kanadensiska ambassaden ?
Var ligger den egyptiska ambassaden ?
Var ligger den finska ambassaden ?
Var ligger den danska ambassaden ?
Var ligger den grekiska ambassaden ?
Var ligger den ungerska ambassaden ?
Var ligger den indiska ambassaden ?
Var ligger den israeliska ambassaden ?
Var ligger den italienska ambassaden ?
Var ligger den nyzeeländska ambassaden ?
Var ligger den norska ambassaden ?
Var ligger den portugisiska ambassaden ?
Var ligger den ryska ambassaden ?
Var ligger den spanska ambassaden ?
Var ligger den nederländska ambassaden ?
Var ligger den turkiska ambassaden ?
Var ligger den brittiska ambassaden ?
Var ligger den amerikanska ambassaden ?
Jag väckte dig .
Detta måste stoppas genast .
Det hände så fort .
Sjutton gastar på död mans kista , yo-ho och en flaska med rom !
Sjutton gastar på död mans kista . - Hej och hå och en flaska med rom !
Succé !
Detta är den femtusende klingonska meningen på Tatoeba !
Vi är hans söner .
Kan du hjälpa mig ?
Jag skrev min första mening på tyska .
Jag föreslog honom att hon skulle bli inbjuden till festen .
Jag skriver en mening på tyska .
Jag försöker översätta .
Jag kan inte leva utan dig .
Jag kan inte se dig .
Jag vet inte varför .
Jag vet inte vad jag vill .
Jag vill lära mig tyska med mina vänner .
Hon talar inte engelska .
Nej , jag är engelsk .
Hans fru är svensk .
Svenska är lätt .
Det är min son .
Min son talar inte svenska .
Jag skriver korta meningar på svenska .
Jag skriver en sång på tyska .
Jag skriver ett brev till min fru .
Jag räknar på tyska .
Jag läser det här brevet .
Algeriet ligger i Nordafrika .
Algeriet är mitt land .
Pfirsichbaeumchen är från Tyskland .
Jag lär mig svenska och tyska .
Du lär dig arabiska .
Var ligger Algeriet ?
Jag vill ha en bok på svenska .
Wenjin är en kinesisk kvinna .
Känner du mig ? – Nej .
Jag misstänkte att han ljög , men det kom inte som en överraskning .
Jag kommer tillbaka om en timme .
Sanningen är att jag älskar dig .
Var bor du ?
Kan du franska ?
Vi ses om två år .
Jag gillar musik , speciellt klassisk sådan .
Jag följer med dig och handlar .
Stranden är ett idealiskt ställe för att barn att leka .
Natten är ju ganska lång , eller hur ?
Stäng dörren när du går .
Fattigdom är ingen skam , men den hjälper ingen fram .
Fattigdom är ingen skam .
Klarar du dig med engelska ?
Tom bor inte här .
Det är någon vid dörren .
Telefonen ringer .
Jag ska studera engelska i eftermiddag .
Patricia kommer att hålla i turneringen .
Livet är vackert .
Jag hatar dig väldigt mycket .
Tom är en mycket stark man .
Vår lärare är alltid i tid till lektionerna .
Jag trodde att jag förstod dig .
Skulle klockan åtta passa ?
Gör gott mot dem som hatar er .
Gören gott mot dem som hata eder .
Bestämt inte .
Tom får rösta .
Hur gick din intervju ?
Jag råder dig att inte åka .
De senaste medicinska framgångarna är anmärkningsvärda .
Det ligger en bok om dans på skrivbordet .
Tom bestämde sig för att läsa juridik .
Jag ska plugga engelska i eftermiddag .
Tom måste välja mellan heder och död .
Jag gör det för att jag måste .
" Varför ska du inte åka ? "
" För att jag inte vill . "
" Skicka mig saltet , tack . "
" Varsågod . "
Det är för mycket att göra .
Jag har huvudvärk .
Ring polisen !
Det ligger inte långt härifrån .
Vi hängde oss alla åt vårt lands utveckling .
Hon kom inte förrän två .
Jag behöver en ny cykel .
Vet du var mina gamla glasögon är ?
Tom skrattade åt Mary .
Det tar oss fem minuter att gå igenom tunneln .
Jag skulle vilja stanna en natt .
När man talar om trollen !
Din cykel är mycket nyare än min .
Var är toaletten ?
Jag studerar på universitetet i Hyogo .
Lektionen börjar inte förrän halv nio .
Vem springer snabbast i din klass ?
Han betonade att tiotusentals människor skulle komma till konserten .
Tom hoppade av sin häst .
Ingen kan undkomma döden .
Jag visade för dem hur man gör .
Min klocka är tio .
Vad betyder det här ordet ?
Det finns många amerikaner som kan tala japanska .
Han spenderade slut på sina pengar .
En ishockeypuck är inte klotformad .
Och inte här heller .
Tom är övertygad .
Jag var väldigt glad .
Jag gillar hundar och min syster gillar katter .
Är du nöjd med resultatet ?
Le nu , gråt senare !
Han tjänar tre gånger så mycket pengar som jag gör .
Jag kan inte hitta Tom .
Har han redan gått ?
Jag ska arbeta under sportlovet .
Är det mig du menar ?
Jag behöver någon för en vuxen .
Saknade du mig ?
Du har köpt fler frimärken än vad som är nödvändigt .
Jag måste gå och handla .
Jag är tillbaka om en timme .
Var är vi ?
Hur mycket förbrukar den här bilen ?
Hela historien är höljd i dunkel .
Jag ska köpa en ny .
Jag kan komma klockan tre .
Han är en bra förlorare .
Jag minns inte hennes namn .
Den paranoida mannen anförtrodde sig inte åt någon alls .
Jag har tappat bort mitt bagage .
Hon var ung och oskyldig .
Jag arbetar här .
Både hans morfar och farfar är döda .
Om det regnar stannar jag hemma .
Där tar du troligen fel .
Tom gjorde det för skojs skull .
Jag trivs verkligen i Georgia .
Hade jag vetat skulle jag ha sagt det till dig .
Skulle jag kunna få använda din telefon ?
Han känner många människor .
Tom förväntade sig inte riktigt att Mary skulle svara på hans fråga .
Det är bara ett talesätt .
Tom bor med Mary i Memphis .
Om hon bara hade vetat att jag var i Tokyo , skulle hon ha hälsat på mig .
Allt är i sin ordning här .
Ursäkta .
Jag skulle vilja hyra en bil .
Hur gick det på din intervju ?
Vi har en reservation klockan halv sju .
Han kom i går för att träffa oss .
Det här är mannen som jag letat efter .
Skulle du vilja dansa med mig ?
Öppna munnen !
Han är redan en man .
Jag vill inte vara rik .
Vem talar jag med ?
Vem pratar jag med ?
New York är en av de största städerna i världen .
Du borde ha avvisat ett sådant orättvist förslag .
Barnuppfostran är en hård uppgift .
Jag känner inte för att äta just nu .
Du kommer läsa det någon annan dag .
Ärligt talat så är hon en opålitlig typ .
Vi satte oss i bilen .
Jag har mycket att göra i dag .
Äter du ofta fisk till middag ?
Nu är det mat !
Varsågod och ta lite tårta .
Kleta inte i bibliotekets böcker .
Drick inte så mycket öl .
Hon hoppade på tåget .
Du borde verkligen inte dricka kranvattnet .
Datorn är en komplicerad maskin .
Hon stod käpprak .
Hon tror alltid på mig .
Har ni några fler frågor ?
Ken vann över mig på schack .
Jag vill ha en båt som kan ta mig långt härifrån .
Jag ville bara kolla min mejl .
" Hon gillar musik . "
" Det gör jag med . "
Skulle jag kunna få tala med fröken Brown ?
Vinden avtog .
Jag var mycket glad .
Sjön ser ut som ett hav .
Jag är vilse .
Kan du hjälpa mig ?
Beskedet kom som en blixt från klar himmel .
Det är regn på väg .
Jag gav dig en bok .
Den gamla gubben ruckar aldrig på sina principer .
Jag trodde att jag sa åt dig att inte komma .
Översätt inte den här meningen !
Vi kunde inte gå med på hans krav .
Hans imponerande tal var som pärlor för svinen .
Jag vill inte gå ut utan jacka en sådan här kall dag .
Prinsessan låg med slutna ögon .
" Tack så mycket " , sa han med ett leende .
Ingen vet om hon älskar flickan eller inte .
Detta är första gången jag ber i en moské .
Det är bäst att du gör det omedelbart .
Jag blir alltid nervös när jag kommer i närheten av henne .
Det är det dummaste som jag någonsin sagt .
Titta på mig när jag pratar med dig !
Hon vill inte prata om det .
Jag märkte det inte förrän i går .
Min tv har slutat fungera .
Jag skulle vilja gå hem nu .
Vad sägs om lite fika ?
Är någon sugen på fika ?
Du står näst på tur för en befordran .
Du är en idiot .
Välj oss !
Kulramen är en kinesisk uppfinning .
Han har en dålig vana att dricka för mycket vin .
Var ligger kaffeaffären ?
Han lyssnade på musik för sig själv .
Nästan alla löv har fallit av .
" Vem är det ? "
" Det är din mor . "
Du ser dum ut .
Han talar franska .
När kommer tåget fram till Yokohama ?
Jag tycker om honom väldigt mycket .
Jag är för gammal för den här världen .
Tom verkar vara en idiot .
Vilken ordbok syftade du på ?
Jag tycker om hundar och min syster tycker om katter .
Jag ser fram emot sommarlovet .
Han kom nyss tillbaka hem .
De darrade som asplöv .
Du kommer inte kunna övertala Tom att göra det där .
Offret låg med ansiktet ned i mattan .
Tom ligger i sängen .
Tom kunde inte tro på det som hänt .
Är det där franska ?
Sånt är livet .
Vänta på er tur .
Jag minns inte hans namn .
Jag älskar det norska språket !
Jag vill inte alls åka .
Han talar inte lika flytande engelska som du .
Varför studerar ni franska ?
Fortsätt bara denna gata framåt ungefär 200 meter .
Jag gick ofta på bio med pappa .
Har ni några syskon ?
De skyndade sig ut ur rummet .
Jag tror att hon är ledig i morgon .
Kan man få byta rum ?
Jag kan inte skylla olyckan på honom .
Du har bättre kondition än jag .
Jag skulle vilja få ett allvarsord med dig .
Tydligen inte .
Hon spenderade slut på sina pengar .
Vilken årstid gillar du mest , våren eller hösten ?
Du borde sova .
Jag trivs verkligen i Georgien .
Det kommer försätta dig i fara .
Katten stirrade intensivt på honom med sina stora , runda , blåa ögon .
Det kommer att bli ganska kyligt .
Han torkade svetten från ansiktet .
Jag lovar .
Han hade få tänder .
Sann kärlek existerar inte .
Varje gång de pratar med varandra blir de osams .
När man talar om trollen så står de i farstun .
Jag har nariga läppar .
Invektiven haglade över honom .
Pojken kikade genom en springa i staketet .
Jag är en pålitlig person .
Pojken är som en miniatyr av sin far .
Hon talar inte lika flytande engelska som du .
I den där affären säljs köksredskap .
Varför läser du franska ?
Hon låg med slutna ögon på soffan .
Han låg med slutna ögon på soffan .
Tom fick slut på bensin .
Vi hyrde en lägenhet .
Hämta mig dagens tidning .
Jag är finsk .
Har jag fått några telefonsamtal ?
Vi träffades under ett ensamt träd .
Han hoppade på tåget .
Det gör inte så ont .
Jag har inte ätit ordentligt på en vecka .
Ingenting .
Strunt samma .
Vem vill ha lite varm choklad ?
Ge mig ett halvt kilo äpplen .
Ingen vill arbeta utomhus under kalla dagar .
Vilka vackra blommor !
Barnet tigger alltid om någonting .
Tom bestämde sig för att skjuta upp beslutet .
Å min sida , hoppas jag att det inte ska regna .
Regnet stod som spön i backen .
Jag vill åka utomlands någon dag .
Han sprang så fort som han kunde .
Titta på skylten framför dig .
Det är inte bra att bryta ett löfte .
Han var tålmodigheten själv .
Jag kan inte leva ett sådant liv .
Vet du vilka färger hon tycker hon ?
Vet du vilka färger han tycker om ?
De snackade hela natten .
Han drunknade nästan i floden .
Hon drunknade nästan i floden .
Jag vill inte ha någon frukt .
Mina ekonomiska bekymmer är över .
Denna byggnad håller på att rasa samman .
Han arbetar på ett laboratorium .
Vet ni hur man öppnar den här lådan ?
Den där klänningen passar dig bra .
Han bor i en lägenhet .
Hon bor i en lägenhet .
Till och med under arbetstid ger jag i lönndom efter för mitt internetberoende .
En hund sprang .
Alla är redo .
Jag tror att han är ledig i morgon .
Varför uppför sig män som apor , och vice versa ?
Jag studerar engelska , eftersom jag ska åka till USA .
Hur tar jag mig till busshållplatsen ?
Du borde slå upp det ordet .
Jag går och klär på mig .
Jag skulle vilja köpa en karta .
Vem stal äpplet ?
Jag missade mitt tillfälle .
Denna fågel lever varken i Japan eller i Kina .
Bättre sent än aldrig .
Hon är min bästa vän .
Vad är bättre än en skål med popcorn och en med glass .
Jag växte upp med att titta på Pokémon .
Schweiz är ett väldigt vackert land och är mycket värt att besöka .
Han blir sällan arg .
Det spelar ingen roll vilket lag som vinner matchen .
Tv : n är på .
Vem tror du att du är ?
Jag fick ett brev från min vän .
Tom behöver köpa en ny regnrock .
Hon är min fru .
Min syster har gett mig en iPhone , men jag vet inte hur man använder den .
Jag missade tåget med bara några minuter .
Är du jänkare ?
Kinesisk filosofi är bäst .
Jag har tappat bort min penna .
Släpp honom !
Låt mig följa dig hem .
Den gamla kvinnan gick upp för trappan med möda .
" Tammi " med två m .
Alltså T-A-M-M-I .
Kan jag få ett kvitto , tack ?
Min pappa tycker om tennis .
Både hennes morfar och farfar är döda .
Bry dig inte om andra .
Det gick ju smärtfritt .
Det är inte mödan värt .
Vem ser efter dina hundar ?
Skynda er .
Annars kommer vi försent till lunchen .
Är det illa ?
Jag är inte färdig än .
Hur var din kväll ?
Du är det vackraste flickan jag någonsin sett .
Det är farligt för dig att simma i den här floden .
Katten är under bordet .
Ärligt talat har jag redan sett den filmen .
Ät upp det där brödet !
Hämta mig en torr handduk .
Glöm inte det .
Jag läser koreanska .
Är du galen ?
Termiter äter trä .
En ishockeypuck är inte sfärisk .
Lyssnar du på mig ?
Han är någonstans i parken .
Han höll på att diska .
Tekniken fallerade och hela tillställningen fick avbrytas .
Han kastade ett öga på sin klocka .
Du är bara en hora .
När farfar pratar om barndomsminnen blir han lätt oratorisk .
Jag ska ta med min son till djurparken i eftermiddag .
De är på god fot med sina grannar .
Har ni några frågor ?
Jag vill förändra världen .
Vänta på din tur .
Av tre hundar är en en hane och två honor .
Hej , Tom !
Bågskytten dödade hjorten .
Om ni vill tala med mig , så ring .
Vi kunde inte gå med på hennes krav .
Vi lyssnar på musik .
Vill du ha mer te ?
Vår skola ligger i den här byn .
Det har aldrig snöat så här mycket .
Ingen vet om han älskar flickan eller inte .
Kragen sitter åt för hårt runt min hals .
Jag kom från Kina .
Jag blir ofta förkyld .
Han tappar alltid bort sitt paraply .
Det här kommer aldrig att ta slut .
De här hörlurarna fungerar inte .
Tom har stor respekt för Mary .
Att vara hemma är inte kul .
Hennes pappa var polis .
Han verkar ha haft ett svårt liv i sin ungdom .
Så blå himlen är !
Men berätta då !
Vi skattade oss lyckliga som överlevde .
Han blir lätt trött .
Tiden är ur led .
Jag tänkte att det var värt ett försök .
Sådant är livet .
Telefonen ringde .
Låt oss hoppas på det bästa i alla fall .
Förutom engelska talar han tyska .
Ingen vet vare sig han älskar henne eller inte .
Hon sa att de var goda vänner till henne .
Har ni något mer att säga ?
Jag säger samma sak om och om igen .
Han väntade på sin tur .
Hon har köpt en ny dator .
Det här är huset , i vilket min farbror bor .
Du är i vägen .
Jag hjälper dig gärna .
Jag vet inte om han är en doktor .
Jag skriver ett brev .
Det skulle jag aldrig ha gissat .
Jag är så upptagen att jag inte kan hjälpa er .
Jag kommer inte ihåg vad hon heter .
Att skriva dagbok hjälper oss att minnas små , dagliga saker .
Titanic krockade i ett isberg .
Hon kommer kanske .
Du kom ändå !
Mamma satt mig i arbete emot min vilja .
Jag trodde att fienden hade dödat Tom .
Tom ligger på backen .
I morgon ska jag åka till Shanghai .
Wikipedia är den bästa encyklopedin på nätet .
Hunden är människans bästa vän .
Vi skyndade oss , så att vi hann med den sista bussen .
Förutom engelska talar hon tyska .
De pratade hela natten .
Jag trodde att jag var trevlig .
Jag beundrade hans generositet .
Jag sparar till en moped .
Hon övertalade honom att göra det fastän hon visste att det inte var en god idé .
Jag ville bara kolla min mail .
Muiriel är 20 nu .
Hur är läget ?
Hur har din dag varit i dag ?
Han vann första pris på schackturneringen .
Mark stöter på allt som rör sig .
Hur säger du det på italienska ?
Vi diskuterade vad vi skulle göra .
Jag vet inte om han är en läkare .
Hon är givmild med sina pengar .
Jag tycker om henne väldigt mycket .
Han är min bästa vän .
Jag vill inte gå till skolan .
Ibland känner jag mig ledsen .
Jag vet att jag kommer att dö .
Det är dig som hon älskar , inte mig .
Jag tycker att du borde vila ; du ser sjuk ut .
Jag var hungrig .
Kan jag använda telefonen ?
Nu kryper vi till kojs .
Engelska och tyska är besläktade språk .
Hon samlar ihop pengar till handpenningen .
Jag sparar till en moppe .
Jag är trött eftersom jag var tvungen att plugga inför ett prov igår natt .
Om du har läst ut boken , så skulle jag vilja låna den .
Han har bott på det där hotellet de fem senaste dagarna .
Hon blev tvungen att förlita sig på sin inre styrka .
Ungefär 9,4 % av jordens yta är täckt av skog .
Hur lång tid tar det till stationen ?
Han du någonsin ätit en bananpaj ?
Han är anklagad för förargelseväckande beteende .
Vad fin det är !
Gjorde du den helt själv ?
Har du läst ut boken ?
Hans kunskaper i kinesiska gjorde att vi kunde genomföra planen smidigt .
Detta är huset där han bor .
Talarens påstående var irrelevant .
Det är ett mycket välbesökt kafé .
Kvinnan hade ett ångerköpt uttryck i ansiktet .
Ett glas kall öl skulle göra gott .
Min bror är bra på tennis .
Hur var din dag ?
Engelska studerar man även i Kina .
Jag är hungrig eftersom jag inte åt frukost .
Det här året erbjuder vi samma språkkurs som i fjol .
Du ser riktigt trött ut .
Ärligt talat så är han en opålitlig typ .
Jag har precis ätit färdig .
Jag gillar inte dina vänner alls .
Han är väl inte här ?
Lämna inte tv : n på !
Jag bad honom om råd .
Jag bad henne om råd .
Dock är det något som överlevandena inte känner till .
Jag ska presentera dig för några vänner som läser tyska .
Det var hans tystnad som gjorde henne arg .
Han har redan gått .
Vad är det du vill säga egentligen ?
Vem uppfanns telefonen av ?
Jag skulle aldrig ha gissat det .
Jag har två äldre syskon .
Han drar ifrån .
Vi ska åka till Estland nästa månad .
Tom ligger på rygg .
De frågade Kate om hon kunde sitta barnvakt åt barnet .
Tom gav Mary en kopp .
Ni borde fråga honom om råd .
Hans pappa var polis .
Talar du italienska ?
Hon kom i går för att träffa oss .
Jag har en hemsk huvudvärk .
Jag tror fortfarande på kärleken .
De gick och fiskade i går .
Var bor din morfar ?
Berätta för mig när han kommer .
Han var tillräckligt dum för att tro det .
Jag skulle vilja att du hjälper mig med en sak .
Påfrestningen börjar ta på henne .
Du ljuger !
I morgon åker han till Kina .
Äntligen lättade molntäcket .
Ni har en telefon .
Ett , två , tre , fyra , fem , sex , sju , åtta , nio , tio .
Vad gör Jon just nu ?
Tom lånade en bok från Mary .
Jag har aldrig sett ett rött kylskåp .
Var det något mer ni skulle få sagt ?
Jag kan inte .
Färgen är lite för mörk .
Det gör ont .
Sluta !
Kolumbus fann Amerika år 1492 .
Detta är Ken .
Han älskar sin hund .
Tom är groggy .
Få bort honom från vägen .
Få bort henne från vägen .
Tom är skild .
Är allt okej ?
Ät det där brödet !
Hon lyssnade på musik för sig själv .
Jag har många blommor .
Några är röda och andra är gula .
Vilket land är störst , Japan eller England ?
Han tror alltid på mig .
Förlåt att jag har orsakat dig så mycket besvär .
De säger att kärleken är blind .
Finns det reserverade platser på tåget ?
Varje år publiceras det många böcker .
Antingen talar vi kinesiska , eller så talar vi inte alls .
Du kanske kommer att lyckas .
Det är molnigare i dag än i går .
Vänta fem minuter , är ni snälla .
Det är inte möjligt !
Det här är den högsta byggnad som jag någonsin har sett .
Hur lång är ni och hur mycket väger ni ?
Vems gitarr är det här ?
Han var allt annat än nöjd med sin egen framgång .
Hur mycket kostar den här radion ?
Fortsätt arbeta .
Du har förändrats .
Det ser värre ut än det är .
Beträd ej gräsmattan !
Oroa dig inte .
Huset är kallt .
Den här fågeln är utrotningshotad .
Jag tar en kopp kaffe , tack .
Elefanter är enorma djur .
Inget är viktigare än medkänsla .
Han kom för att träffa oss i går .
Hon kom för att träffa oss i går .
Jag skulle gärna resa världen runt .
Jag tror att jag ska stanna här .
Du dricker för mycket kaffe .
Jag skulle vilja veta anledningen .
Han bor hos sina föräldrar .
Han var på väg till skolan .
Hon skrattar sällan , om ens någonsin .
Tom är inte en lat pojke .
I själva verket arbetar han hårt .
Han kan inte kontrollera sina känslor .
Hon kan inte kontrollera sina känslor .
Han försökte att studera hela natten , dock i onödan .
Varför gjorde han det där ?
Varför gjorde han så ?
Jag trodde att han var sjuk .
Jag jobbar här .
Dörren går inte att stänga .
Det här problemet är svårlöst .
Vi visade honom bilder från Alperna .
Du är människa .
Du är en människa .
Du ser verkligen trött ut .
Ingen vet om han älskar henne eller inte .
Mor köpte två flaskor apelsinjuice .
När åkte du till Rom ?
Trots att det regnade så spelade vi fotboll .
Vi var på bio i går .
Skolan är tråkig .
Romanerna han skrev är intressanta .
Någon har stulit alla mina pengar .
Jag hade tur .
Han är givmild med sina pengar .
Det var fler än en som blev uppbragta över politikerns skamlösa skattesmitning .
Har hunden fått vara ute någonting då ?
De får veckolön .
Jag ger dig mitt ord .
Vart går du oftast och klipper dig ?
Jag föredrar komedier framför tragedier .
Vilken av dessa hundar är din ?
Skicka saltet .
Det är inte lätt att lösa problemet .
Var bor din farfar ?
Tom hade tur som hittade sina nycklar .
Det är min fru .
Det är för varmt .
Sophies finger blödde så mycket att blodet droppade ner på marken .
Jag är väldigt känslig emot kyla .
Skulle jag kunna få ett till täcke ?
Jag har varit upptagen hela dagen .
Du kan lita på Jack .
Jag studerar spanska den här terminen .
" Nyckeln sitter i låset " , tillade mannen .
Jag behöver pengar .
Vi gick för att simma i floden .
Var inte rädd .
Jag fick nästan full poäng .
Han höll sitt löfte .
Det här läkemedlet passar inte mig .
Den här medicinen passar inte mig .
Vissa tycker att hemlagat är nyttigare än restaurangmat .
Han hade inte ätit på två dagar .
Jag fick en skriftlig inbjudan .
Jag har några engelskspråkiga böcker .
Han var så hungrig att han åt tallriken tom utan en sekunds tvekan .
De kunde bara lyssna .
Detta är mannen vars resväska jag fann .
Du behöver inte stressa med att byta kläder .
Vi har nämligen ingen anledning att skynda oss .
Min fru är läkare .
De lyssnar inte alltid på sina föräldrar .
De lyder inte alltid sina föräldrar .
Jag vill inte bli utnyttjad .
Du kan välja vilken bok du vill .
Ni får välja vilken bok som helst .
Jag hittade ett väldigt trevligt ställe i går .
Det tjänar inte att fastna i gamla spår .
Tåget stannar på varje station .
Skulle jag kunna få mer potatismos .
Han ville gå hem , men gick vilse på vägen .
Nu är det officiellt .
Jag ska åka till Paris i höst .
När man har feber är det bäst att stanna hemma .
Vi tycker inte om regn .
Han åkte till Tokyo i går .
Jag åkte till London .
De diskuterade problemet .
Vi ses vid huset !
Skulle herr Virtanen vilja ha lite kaffe ?
Jag kan fortfarande inte bestämma mig om jag ska åka dit eller inte .
I morgon ska jag visa dig biblioteket .
I ' ll show you the library tomorrow .
Han ser ut som en ärlig person .
Skulle du kunna hjälpa mig en sekund ?
Han påminner särskilt om sin mor .
Hon påminner särskilt om sin mor .
Han är ett huvud längre än jag .
Hon är ett huvud längre än jag .
Hon är ett huvud längre än mig .
Han är ett huvud längre än mig .
Hur mycket kostar trästolen ?
Jack samlar på frimärken .
Han förstår Er inte .
Hon förstår Er inte .
Jag ser en man mellan träden .
Finns den här i blått ?
Hur var vädret i går ?
Hurdant väder var det i går ?
Jag förstår inte det där ordet .
Det där ordet förstår jag inte .
Vad vill du äta till lunch ?
Jag tycker inte om hundar .
Jag tycker inte om eldig mat .
Jag tycker inte om stark mat .
Fråga Alex .
Sådan här musik är inte min grej .
Gör det genast , så att du inte glömmer .
Tom vilar .
Vi är båda studenter .
Jag har ingen vodka .
Jag har inte tid att läsa .
Vi röstade emot förslaget .
Katter ser i mörker .
Just då stannade bussen .
Jag minns inte hans förklaring .
Vems cykel är det där ?
Han ögon är blåa .
Han har redan ätit .
Hon har redan ätit .
Jag vill inte vänta så länge .
Vi åker när det slutat regna .
När man är hungrig smakar allting gott .
Kom hit .
Det är farligt att bada i den här floden .
Bort med armbågarna från bordet .
Varför köpte du en så dyr ordbok ?
En kanin springer i trädgården .
Jag är på balkongen .
Den här klockan är mycket bättre än den där .
Jag råkade glömma telefonladdaren hemma .
Problemet med den svenska animationsbranschen är att den i stort sett är icke-existerande .
Tror du att vi borde överge skeppet ?
Jag har precis kommit hem .
Min far är på promenad i parken .
Hon säger att hon inte dejtar någon just nu , men jag tror inte på henne .
Tom dricker inte öl hemma .
Om en dörrvakt bär ditt bagage , glöm inte att ge honom dricks .
De simmade .
Vi drack en hel del .
Vi drack mycket .
Vad är det för fel på dig ?
Känner du någon som var på det där skeppet som sjönk ?
Skeppet var inte redo för strid .
Var är kaptenen för det här skeppet ?
Varför är du inte redan ombord på skeppet ?
Jag kände att jag bara var tvungen att komma av skeppet .
Du blev tillsagd att stanna på skeppet .
Det här är det bästa skepp som jag någonsin varit på .
Tom tittade ut genom fönstret på skeppet som kom in i hamnen .
Det är ingen på det här skeppet förutom oss .
Hur många människor var ombord på det där skeppet ?
Är Tom fortfarande kapten över ditt skepp ?
Tom föddes på ett skepp .
Vem är kapten över det här skeppet ?
Vem är kapten över detta skepp ?
Skeppet har inte ens dockat än .
De såg antagligen vårt skepp komma in i hamnen .
Tom sa att han läste en bok om det här skeppet .
Jag minns att jag var på ett skepp när jag var bara fem år gammal .
Hur långt borta tror du att det där skeppet är ?
Skeppet genomsöktes noggrant , men inga illegala droger hittades .
När ska skeppet anlända ?
När ska skeppet komma fram ?
Jag har rätt att vara på det här skeppet .
Vi går tillbaka till skeppet .
Vi måste gå tillbaka till skeppet .
Vårt skepp blev inte skadat i striden .
Jag undrar vart det där skeppet är på väg .
Var kom det där skeppet ifrån ?
Vi ses igen när vi är tillbaka på skeppet .
Skeppet börjar sakta att röra på sig .
Det här är en bild på skeppet som jag var på .
Tom berättade för oss att det var ett gammalt skepp .
Vi kommer att söka genom hela skeppet .
Vi ska söka genom hela skeppet .
Jag kan köpa en bil med de här pengarna .
Mayuko har inte sovit tillräckligt .
Hän bestämde sig för att inte gå på festen .
Som tur är har jag tillgång till ett enastående bibliotek .
Hans nya teori är utom mitt förstånd .
Jag kan inte förstå hans nya teori .
Jag började inse , att jag hade missförstått honom .
Jag tycker inte om att tala inför människor .
De tillbringade en underbar tid tillsammans .
De hade det underbart tillsammans .
Hon är äldre än honom .
Vad tittar du på ?
Ska det regna i morgon ?
Hon blandar ofta ihop socker och salt .
Hon var förkyld och nös ideligen .
Fågelkvittret hördes lång väg .
De nykläckta fågelungarna var alldeles duniga .
Fågelungarna hoppas omkring i buren och flaxade intensivt med vingarna .
Katten stirrade med stor intensitet på när fågelmamman matade sina ungar .
Den brunmaskade kattungen kröp försiktigt ned i bädden bredvid den stora , svarta labradorhanen .
Hennes självsvåldiga beteende möter ofta kritik i samarbetskrävande situationer .
De självutnämnda proffsen var mer eller mindre initierade i företeelsen .
Månne inte snön smälter snart .
Månne bensinpriset skjuter i höjden i sommar .
Kan han månne ha ett slaviskt språk som modersmål ?
Barnet blev tvunget att förlika sig med det faktum att mamma bestämmer .
Han gjorde ett tappert försök att förkväva de känslor som kokade inom honom .
Han har svårt att se framtiden med tillförsikt .
Han har ingen positiv syn på framtiden .
Vi hade stora svårigheter att hitta busshållplatsen .
Den livslust varmed hon bekämpade sjukdomen var beundransvärd .
Det skramlade till av mynt som slog emot varandra i hennes ficka .
Kulen , gråkall , råkall , kylig , ruskig och ruggig är alla synonyma ord för ett väldigt otrevligt väderförhållande .
De fick låna påslakan .
Han slog på spisen och satte ungen på 200 grader .
Spisplattan var fortfarande varm efter en kvart .
Hon blev tacklad och föll till marken .
Barnpassning kan vara ytterst tålamodsprövande .
Då får det vara .
Han är en mycket fåordig man .
De stod med böjda knän och tittade på marken .
Han fick ett undvikande svar .
Barnen dök i bassängen .
Det gläder mig att höra hur bra det går för dig !
Det är om något ett glädjeämne .
Den här åkattraktionen är parkens riktiga dragplåster .
Det halkade bara ur mig !
Stereon dunkade på högsta volym .
Varför läser jag isländska ?
Varför studerar jag isländska ?
Varför lär jag mig isländska ?
Grytan stod och puttrade på spisen .
Jag ska skjuta honom .
Jag tror jag ska gå och lägga mig .
Det är dags att inse att det är omöjligt .
Vi kommer aldrig att klara det .
Jag vill inte tillbaka .
Dörrar är inte så illa som du tror .
Dörrar är inte så dåliga som du tror .
Särskrivning är en allt för vanlig företeelse i det svenska språket .
Jag känner mig småfrusen .
Jag försade mig .
Hon glömde paraplyt hemma och blev helt genomblöt i regnet .
Han blev halvt ihjälslagen .
Han blev slagen blodig .
Sluta mucka gräl nu !
Generellt sett lever kvinnor längre än män .
En vän i handen är bättre än tio i skogen !
Kan du skicka mig den där grunkamojen ?
Jag såg du-vet-vem i dag på torget .
Jag ska precis till att skriva en mening på tyska .
Jag kommer att skriva en mening på tyska .
Jag ska skriva en mening på tyska .
Om ett mänskligt liv är konvext , kan vi optimera det .
Hon nekade mitt önskemål .
Den här jakten är väldigt dyr .
Den här yachten är väldigt dyr .
Denna lustjakt är väldigt dyr .
Hon har möjligheten att arbeta !
Han har möjligheten att arbeta !
När jag fantaserade fram fantasibilder fantaserade jag att min fantasiförmåga fantaserade alla bilderna .
Tänk dig att ens fantasiförmåga fantaserar fram fantasier som man inte ens kan fantasera om .
Confucius sade : " Den som inte dricker te är en dåre . "
Jag hittade en mycket intressant hemsida som lägger fram fullständiga texter om isländska sagor , av vilka några också är översatta till engelska och danska .
Jag skickade ett brev till Steina på isländska .
De vill att vi ska tro att vi lever i en demokrati .
Vad ska du göra på Halloween ?
Kriget tog slut 1954 .
Jag gillar tecknat .
Jag gillar serieböcker .
Jag gillar manga .
Tranan kikade på tranornas halsar .
Tranan kikade på tranornas gurkor .
Det är enkelt att göra och det är billigt .
Jag gör det här för hennes skull .
Är du redo för Halloween ?
Om det inte låter engelskt är det inte engelska .
Det jag skrev är inte engelska .
Jag ska göra mitt bästa .
Låt inte den här informationen läcka ut .
Var är min tidning ?
Vi blev tillsagda att stanna på skeppet .
Tom är arg .
Sötningsmedel har till mångt och mycket samma effekt som socker .
Vår lärare sa till oss att vi bör göra vårt bästa .
Jag undrar vem som namngav detta skepp .
Jag är kapten över detta skepp .
Vilket skepp kommer du med ?
Vilket skepp kom Tom med ?
Deras skepp ligger fortfarande i hamn .
Kom prick klockan tio .
Jorden är mindre än solen .
Tom kan inte sitta i bilen längre än tio minuter innan han blir åksjuk .
Jag fick sendrag i vänstra benet .
Han reste utomlands på statens bekostnad .
Blodet stelnade i ådrorna på honom .
Något liknande hände mig förra året .
Han tog sin tid .
Orkanen Sandy är på väg .
Skulle du kunna vara tyst , tack ?
Vi försökte att kontakta det andra skeppet .
Skoldagen kändes som en evighet .
Det där släktdraget går i rätt nedstigande led .
Den stökiga eleven blev utskälld efter noter .
Det slog mig att du kanske inte heller har sett den filmen .
Han föreställer sig allt möjligt .
Vi fann böckerna slängda huller om buller på golvet .
Hon fick en futtig summa i ersättning för skadan .
De accepterar inga avvikelser från mönstret .
Han avlägsnade sig från platsen .
Flickan skriver dagbok i hemlighet .
Skeppet kapsejsade .
Jag rörde ingenting .
Fienden förstörde många av våra skepp .
Varför är du på det här skeppet ?
Var är skeppet nu ?
Jag behöver de här pengarna .
Jag behöver dessa pengar .
Bredvid järnvägsstationen ligger ett solrosfält .
Hur många gånger ska jag behöva berätta för dig att du inte får skrika här inne ?
De har sagt upp sitt telefonabonnemang .
Jag vill egentligen bara skaffa vänner .
Jag arbetade ihjäl mig i det där projektet .
Är det något särskilt som du vill ha att dricka ?
Är det något särskilt som du vill ha att äta ?
Är det något särskilt som du vill titta på ?
Är det något särskilt som du vill höra ?
Är det något särskilt som du vill ?
Är det något särskilt ?
Livet är för kort för att lära sig tyska .
Det är mycket vatten i dammen i dag .
Förut gick jag varje dag på morgonpromenad .
Jag tycker om att resa .
Vad du vad han sa ?
Pratar du med din hund ?
Älskar du honom fortfarande ?
Älskar du henne fortfarande ?
Han älskar henne fortfarande .
Han älskar honom fortfarande .
Hon älskar henne fortfarande .
Hon älskar honom fortfarande .
Det finns goda grunder för att tro på vad han säger .
Vi kallar vår hund för Johnny .
Vår hund kallas för Johnny .
När gifte du dig ?
Varför är hon så olycklig ?
Av vilken anledning är hon så olycklig ?
Jag använder datorn .
Jag använder dator .
Jag använder en dator .
" Är du lärare ? "
" Ja ! "
För länge , länge sedan levde det på en liten ö en gammal kung .
När slutar din lektion ?
Kan du tala kinesiska ?
Kan du prata kinesiska ?
Kan du kinesiska ?
Det här är ett trähus .
Detta är ett trähus .
Jag skulle vilja ha kaffe .
Nu när jag tänker på saken så levde vår familj ett mycket eländigt liv .
Vare sig den är vit eller svart så är en katt som fångar möss en bra katt .
Jag måste få ordning i skallen .
Jag måste samla mina tankar .
Jag måste reda ut mina tankar .
Jag fryser .
Om jag var du skulle jag inte bry mig om det .
Är det svårt att prata engelska ?
Är det svårt att tala engelska ?
Tänker du ofta tillbaka på din barndom ?
Varje dag cyklar jag eller tar bussen till jobbet .
Vem är han ?
Hans rum var i oordning .
Mike är inte bra på baseboll .
Mike är dålig på baseboll .
Stäng av tv : n .
Det här kaffet smakar diskvatten .
Håll käften och lyssna , unge .
Jag tänker bara på dig .
Du måste ta med dig ditt pass till banken .
Du ser uttråkad ut .
Om jag var du skulle jag följa hans råd .
Jag är en realistisk person .
Det kan hända att han inte kommer .
Det kan hända att hon inte kommer .
Han kanske inte kommer .
När jag var ung , var jag tvungen att arbeta hårt .
Jag hade hans namn på tungan , men fick inte fram det .
Han måste ta hand om sin mor .
Hon måste ta hand om sin mor .
Läs av mätaren .
Jag råkade glömma att låsa förrådet .
Efter en hetsig diskussion gjordes en kompromiss .
Rökarna får i framtiden röka i rökhörnan .
Jag lärde mig det av dig .
Var snäll och ge mig lite mer kaffe .
Skulle du kunna förklara vad det här är ?
Klassisk musik är inte min grej .
Mormors gamla armbandsur har legat och skräpat i byrån i åratal .
Vem skrev den här dikten ?
Vi försökte kompromissa med dem .
Om min bror vore här , skulle han veta hur man gör .
Du har för vana att överdriva allting .
Du har en vana att överdriva allting .
Lägg allt i min korg .
De lade stor uppmärksamhet vid hans ord .
Han är bra på franska , men mycket bättre på engelska .
Det skrivs lika på båda språk .
Det skrivs lika på båda språken .
Han är rik , men desto viktigare : han är väluppfostrad .
Han stal mina pengar från förvaret .
Hon stal mina pengar från förvaret .
Alla hennes pengar stals .
Alla hans pengar stals .
Hon slank ned pengarna i min ficka .
Han slank ned pengarna i min ficka .
Hon smällde igen dörren .
Han smällde igen dörren .
Hon slängde igen dörren .
Han slängde igen dörren .
Kan ni ringa igen senare ?
Okej , men bara på ett villkor .
Kanske någon annan gång .
De åt currykyckling till middag .
Kylan bildade snökristaller på fönstren .
Det finns ingenting värre än telefonförsäljare .
Han lutade sig tillbaka i fotöljen och läste en bok .
Hur kommer det sig att du inte berättar detta förrän nu ?
Jag kan tyvärr inte komma förrän i morgon .
Kommer de redan ?
Sluta skälla !
Alla tavlor i rummet hängde på sned .
Hon är helt utom sig av iver .
Mörkret faller tidigt den här tiden på året .
I skymning är det stor chans att få se vilda djur .
Viltstängsel hindrar viltolyckor .
Viltolyckor är vanliga när det är mörkt och halt ute .
Vägföret är inte det bästa , men vi måste ge oss ut ändå .
Är vi framme snart ?
Rattfyllerister ligger ofta och kör uti väggrenen eller nära mittstrecket .
Den gamle mannen berättade att andra bilister hade tutat på honom i rondellen , och de yngre släktingarna förstod genast att han både kört långsamt och i fel körriktning .
Glöm inte att dra i handbromsen .
Lägg ur växeln och rulla .
Är ni inte trötta ?
Är ni inte trött ?
En japansk trädgård har vanligtvis en damm .
En bra mening är bättre än två dåliga .
Hur lång ledighet kommer du att ha i jul ?
Hur länge kommer du att vara ledig i jul ?
Jag litar mer på en tjuv än på honom .
Det finns faktiskt ingenting som du kan göra åt saken .
Jag varnade honom för faran .
Hon sa själv att hon inte skulle bli kär i någon igen .
Min mor nynnade för sig själv medan hon stökade på med matlagningen i köken .
Jag tog hans närvaro för givet .
Jag gav dem ett tusen yen var .
Jag kan inte göra det ogjort .
Någon tappade sin plånbok .
Någon tappade en plånbok .
Genast lämnade fåglarna sina bon .
Flygplanet lyfte för tio minuter sedan .
Vilken tunnelbanelinje går till stadskärnan ?
Vilken tunnelbanelinje går till centrum ?
Rock tilltalar unga män och kvinnor .
Tom har för mycket arbete att göra .
Britterna trodde att amerikanerna överträdde deras lag .
Britterna tyckte att amerikanerna överträdde deras lag .
Har Jane lämnat Japan för gott ?
Har du tappat vettet ?
Hon betalade för att gå på konserten .
Jag skriver en roman .
Om han inte går i skolan tänker jag inte prata med honom längre .
Läraren tolkade meningen åt oss .
Ge mig en av dina bilder , tack .
Han slutade aldrig att skriva .
Jag antar att vi borde gå nu .
Vi försöker .
Det är första gången jag parkerar min bil i skogen .
Jag älskar naturen , men jag avskyr insekter .
Kan du inte tala engelska ?
Han gick ut i regnet .
Jag är gift och har två barn .
Hur såg rånaren ut ?
Jag tror inte att din teori håller .
Vad skrev du igår ?
Han satt i stolen .
De fortsatte att prata , till och med efter att läraren kom in .
Det här är Ken .
Han älskar sin hund .
Rita ett streck på ditt papper .
Ge mig ett exempel till .
Rör er inte !
Al Smiths föräldrar kom från Irland .
Detta används fortfarande dagligen .
Hon började springa .
Tom arbetar inte lika hårt som han brukade .
De försökte fly .
Jag ska strax gå .
Vill du göra mig sällskap ?
Jag lade på och ringde henne igen .
När jag frågade honom efteråt verkade det som han inte hade menat det som ett skämt .
Och till råga på allt fick jag sparken .
Han deltog i en nätundersökning .
Hon valde skorna som passar till klänningen .
Hon valde skorna som matchar klänningen .
Nu har de skickat datorn .
Det här är ganska exakt .
De är oss på spåren !
Vi klagar alltid .
Det där är faktiskt riktigt elakt .
Vad vill du berätta för oss ?
Vad vill du titta på ?
Var är resten av pengarna ?
Vad hände med resten av maten ?
Jag trodde Tom vad en fullständig idiot .
Vi kan inte bevisa att Tom ljuger , men vi är ganska säkra på att han gör det .
Tom ljuger .
Jag gjorde inte det som han sa att jag gjorde .
Det är tydligt att någon ljuger .
Jag undrar vem av er som ljuger .
Tom ligger på en stor sten .
Varför tar du på min flickvän ?
Varför rör du min flickvän ?
Vad vill du ska hända ?
Vad vill du att jag ska göra ?
Jag ville bara prata med Tom .
Jag väger bara 45 kilo .
Jag var bara där en gång .
Jag gick bara dit en gång .
Jag önskar bara att jag kunde vara så lycklig som du verkar .
Jag önskar bara att jag kunde hjälpa er alla .
Om det bara var så enkelt .
Jag önskar bara att det var så enkelt .
Jag önskar bara hjälpa .
Jag vill bara vara till hjälp .
Jag önskar bara att Tom vore här .
Jag önskar bara att Tom kunde vara här .
Om det bara vore så enkelt .
Jag struntar hellre i skolan och spelar tv-spel istället .
Tamy upptäckte ett misstag i meningsbyggnaden .
Jag är så bråttom att jag inte kan hjälpa Er .
Jag är så upptaget att jag inte kan hjälpa Er .
Skulle jag kunna få lite mer mjölk i kaffet , tack .
Han är ingen poet , men en författare .
Skulle ni vara så snäll och öppna dörren åt mig ?
Skulle du vara så snäll och öppna dörren åt mig ?
Hon avbröt oss när vi höll på att prata .
Han avbröt oss medan vi pratade .
Han gillar att lyssna på radio .
Det är alldeles rimligt .
Farfar började bli gammal , så han pensionerade sig .
Farfar började bli gammal , så han gick i pension .
Farfar har blivit till åren .
Stig på bussen en och en .
Han var mer än kung .
Jag hoppas att jag blir sångare .
Ett egendomligt ljud fick honom att kliva ur sängen .
Ett egendomligt ljud fick henne att kliva ur sängen .
Jag hoppas att det blir en sångare av mig .
Det är min väska .
Under förra året skedde det många trafikolyckor .
Kärleken till konsten förde honom utomlands .
Det här är min väska .
Det där är flickan som jag känner väl .
Jag antar att du är beredd att ta risken .
Jag fick ett brev som underrättade mig om hans ankomst .
Hon skrek till av förvåning .
Du behöver inte prata så högt .
Det finns ingen anledning att prata så högt .
Trots att de släppte datorn från fjärde våningen så gick den inte sönder .
Hör du mig ?
Hur ser du om någon är en löpare ?
Hur vet du om någon är en löpare ?
Varför denna uppståndelse ?
Varför detta tumult ?
Varför detta ståhej ?
Varför detta rabalder ?
Det var ett himla kackalorum där inne !
Han hann , men hon hann inte .
Jag fick min välförtjänta lön .
Han skyndade sig in i bilen .
Han dröjde här en stund .
Han stannade här en stund .
Han var kvar här en stund .
Varför dröjde du så länge ?
Jag försöker igen .
Lunchen är klar !
Middagen är klar !
Middagen är färdig !
Tyngd av blötsnö rasade altantaket till slut in .
Vart anger riktning och var anger position .
Var är han ?
Vart går han ?
På flygplatsen fanns hundratals taxibilar , alla på jakt efter kunder .
Skulle du vilja göra mig sällskap på en promenad i parken ?
Han är en god simmare .
Hon är en god simmare .
Hon simmar väldigt bra .
Sätt på tv : n .
Går det bra om jag sätter på tv : n ?
Går det bra att jag sätter på tv : n ?
Stör det dig om jag sätter på tv : n ?
Skulle du kunna sätta på tv : n ?
Jag satt och tittade på tv när jag råkade somna .
När jag tittar på tv blir jag genast sömnig .
Tigern rymde från djurparken .
Enligt min klocka så är hon fyra nu .
Ska vi träffas i morgon ?
Jag känner din bror väl .
Jag kom hit i går .
Försöker du stöta på mig ?
Folk som har varit med om så kallade ' lucida drömmar ' beskriver dem ofta som ' verkligare än verkligheten ' .
De beskriver också verkligheten efter att de vaknat från en ' lucid dröm ' som ' en nyckfull dröm ' .
En av tigrarna rymde från djurparken .
En av tigrarna rymde från zoot .
Han måste komma söderifrån .
Många tror att fladdermöss är fåglar ..
Många människor tror att fladdermöss är fåglar .
Marys meningar är lätta att översätta .
En tiger har rymt från zoot .
En tiger har rymt från djurparken .
Hon går sällan ut .
Hon vill ha en fjärde generationens iPad .
Kan du simma lika snabbt som han ?
Eleverna lyssnar på en historieföreläsning .
Den här stolen är ful .
Tom är inte den gitarrist som han brukade vara .
Orkidén trivs bäst om den får stå i fönstret .
De erbjöd gästerna lite kaffe .
Tom stängde av tv : n .
Tom kan bara inte komma överens med Mary .
Grönt står för hopp .
Jag har läst engelska i fyra år .
Jag har studerat engelska i fyra år .
Jag står inte ut med det här oljudet längre .
Wenjin är kinesiska .
Hon är en ängel .
Jag har inte läst boken och inte vill jag göra det heller .
Här är en mening , med stavelseantalet , som i en haiku .
En trappa och en trapp är nästan samma sak .
Den förstnämnda finns utomhus och den sistnämnda inomhus .
I Sundsvall kallas trappa för bro .
De flesta människor som äter med gaffel lever i Europa , Nordamerika och Sydamerika ; människorna som äter med pinnar bor i Afrika , Mellanöstern , Indonesien och Indien .
Jag gick till fots .
Det är mycket farligt att gå här om nätterna .
Din bror ber om hjälp .
Skriv din dagliga rapport i dag .
Landet har gemensamma gränser med två andra länder .
Jag försökte , men jag misslyckades .
Dessa blommor blommar tidigare än andra .
Våg efter våg rullade upp på stranden .
Våg efter våg böljade in på stranden .
De säljer diverse varor i den affären .
Valresultatet kommer snart att analyseras .
Jag behöver en blyertspenna .
Jag kan låna en av dina ?
Jag behöver en blyertspenna .
Kan jag låna en av dina pennor ?
Jag skulle vilja träffa dig igen nästa vecka .
Det är en katt i köket .
Det finns en katt i köket .
Talar han franska ?
Talar hon franska ?
Pratar han franska ?
Pratar hon franska ?
Han sa att han hade mycket pengar .
Hon sa att hon hade mycket pengar .
Under många år vände han på vartenda öre för att kunna spara pengar .
Hon jobbade flitigt för att kunna tjäna mycket pengar .
Det är dags att gå och lägg sig .
Jag är italiensk .
Jag har inte ens råd att köpa en begagnad bil .
Affären är öppen hela dagen .
Grekiska är inget enkelt språk .
Grekiska är inget lätt språk .
Han är ung , men han måste försörja en stor familj .
Hon är ung , men hon måste försörja en stor familj .
Till en början förstod jag inte varför .
Hunden är hemma .
Jag blir alltid förkyld om vintrarna .
Han är den sista som skulle prata illa om andra .
Hon är den sista som skulle prata illa om andra .
Jag har aldrig hört talas om den här skådespelaren .
Jag lovar .
Jag kommer aldrig att göra det igen .
Jag föredrar cola framför kaffe .
Finns det mjölk ?
Har du någonsin snarkat ?
Vad lång Tony är !
Vilken lång grabb Toni är !
Kom strax tillbaka .
Kom snart tillbaka .
Du släcker väl ljuset när du lämnar rummet ?
Det som han sa hände , det hände .
Så snabbt som möjligt .
Yumi talar riktigt bra engelska .
Han hoppade över diket .
Hon hoppade över diket .
Han sa att jag skulle kunna använda hans rum .
Hon sa att jag skulle kunna använda hennes rum .
Tom slutade att röka .
Hon börjar bli gammal .
Hon har blivit gammal .
Du borde läsa en sådan bok som han läser just nu .
Ingen tror på vad jag sa .
Ingen tror på vad jag säger .
Han frågade mig om jag ville åka utomlands .
Nej , jag tittar inte på CNN .
Var ligger damernas ?
Jag har mitt eget sovrum hemma .
Skriv endast ut jämna sidor , tack .
Det finns femtio stater i Amerika .
Amerika har femtio stater .
Han betedde sig som ett barn .
Jag trodde att Tom skulle sova över i Boston .
Jag trodde att Tom skulle stanna lite längre .
Jag trodde att Tom skulle tala bättre franska än Mary .
Jag trodde att Tom skulle sova till mitt på dagen .
Jag trodde att Tom skulle komma .
Jag trodde att Tom skulle dyka upp .
Jag trodde att Tom skulle säga det .
Jag trodde att Tom skulle säga hej .
Jag trodde att Tom skulle säga hej till Mary .
Jag trodde att Tom skulle komma ihåg .
Jag trodde att Tom skulle minnas .
Jag trodde att Tom skulle plantera de där blommorna nära eken .
Jag trodde att Tom skulle få panik .
Jag trodde att Tom skulle gripas av panik .
Jag trodde att Tom skulle råka i panik .
Jag trodde att Tom skulle bli panikslagen .
Jag trodde aldrig att Tom skulle sluta prata .
Jag trodde aldrig att Tom skulle hålla käften .
Tack så mycket för att ni bjöd in mig .
Tack så mycket för att du bjöd in mig .
Det är dödligt gift !
Du får inte röra vid konstverken .
Du får inte vidröra konstverken .
Du får inte röra konstverken .
Jag tittade på tv i morse .
Skulle du bara kunna berätta för herr Tate att Helen har kommit för att träffa honom .
Vintertidtabellen har trätt i kraft .
Vintertidtabellen har börjat gälla .
Ring mig i morgon .
Han petar sig i näsan .
Hon petar sig i näsan .
Jag har precis flyttat .
Ljug inte !
Dockan stod i hörnet av rummet , täckt av damm .
Han har tio barn .
Hon har tio barn .
Jag dekorerar gärna mitt rum med blommor .
Tom dök aldrig upp på jobbet i dag .
Tom dök aldrig upp på arbetet i dag .
Säg Mexiko och tankar går till tacos .
För länge sedan fanns här en bra .
För en lång tid sedan fanns här en bro .
Jag känner inte den här staden så väl .
Jag känner inte till den här staden så väl .
Tycker du om den här staden ?
Isen var så tjock att jag kunde gå på den .
Tom arbetar på naturskyddsverket .
Tom arbetar på miljöskyddsnämnden .
Tom arbetar på miljöskyddsstyrelsen .
Tom arbetar på miljövårdsmyndigheten .
I dag har jag fruktansvärt mycket läxor .
Om det inte finns någon lösning , så finns det inte heller något problem .
Finns det ingen lösning , finns det inget problem .
Ha alltid en hink vatten till hands , i händelse av en brand .
Musik är hennes passion .
Musik är hans passion .
Vi kunde inte följa hans logik .
Jag tackar för inbjudan .
Det där kan inte vara bra för din hälsa , inte sant ?
Det där kan inte vara bra för hälsan , inte sant ?
Vet du vad hon heter ?
Vad du vad han heter ?
Vi män har vant oss att vänta på kvinnorna .
" Min pappa dricker inte sake . "
" Inte min heller . "
Maria hatar sitt jobb av många anledningar .
Maria hatar sitt arbete av många anledningar .
Thomas tittar på film .
Det kan hända att han inte kommer att lyckas .
Det kan hända att hon inte kommer att lyckas .
Det är en påfågel på gården .
Det står en påfågel på gården .
Han är ett krigsbarn .
Jag är inte intresserad av modern konst .
Den som inte älskar sig själv kan inte heller älska andra .
Tack , allt är bra där .
Hon har inte sett honom på länge .
Om du har följt vad jag har skrivit tidigare .
Jag lämnar tillbaka boken så fort jag kan .
Hon har inte råd med det .
Jag måste sova .
Detta är hans enda chans .
Detta är hans enda möjlighet .
Jag skulle vilja öppna ett checkkonto .
Den här bilen går på alkohol .
Under soffan finns många dammråttor .
Det finns många dammråttor under soffan .
Vilka skolor härstammar från det Buddistiska tänkandet ?
Jag har en flickvän .
Jag blev Toms vän .
Jag fick just en vän .
Jag kanske är din enda vän .
Jag önskar att jag hade fler vänner .
Jag har en vän vid namn Tom .
Jag har en vän vars namn är Tom .
Jag har en vän som heter Tom .
Jag sov inte bra i natt , så jag har inte så mycket energi i dag .
Mina planer misslyckades rejält .
Regeringens politik misslyckades kapitalt .
Mina planer misslyckades kapitalt .
Alla har rätt till sin egen åsikt .
Men ibland är det bättre att hålla den för sig själv .
Tom är en av mina vänner .
Tom är en av mina närmsta vänner .
Jag är Toms vän .
Jag saknar mina vänner .
Jag är Marys pojkvän .
Jag var tillsammans med vänner hela förra natten .
Vem är det som läser ?
Kan jag få se på menyn ?
Skulle jag kunna få ett par ostsmörgåsar ?
Skulle jag kunna få ett glas mjölk , tack ?
Skulle jag kunna få ett glas öl , tack ?
Skulle jag kunna få ett glas vin , tack ?
Jag skulle vilja köpa några vykort .
Det är en buss här .
Det är en krona här .
Det är en smörgås här .
Det finns en busshållplats här .
Det är ett par här .
Det finns ett par här .
Det står ett glas här .
Det finns ett vykort här .
Det finns ett glas här .
Det finns ett hotell här .
Skulle du kunna kolla vad som går på bio nästa lördag ?
Hon klär sig alltid i svart .
Han klär sig alltid i svart .
Hon bär alltid svarta kläder .
Han bär alltid svarta kläder .
Jag uppfattade inte riktigt ditt ärende .
Jag säger det till dig för sjuttioelfte gången – Nej !
Tokyo , som är Japans största stad , är vaken tjugofyrasju .
Har ni någon arbetslivserfarenhet ?
Han tappade bilnyckeln .
Röker ni ?
I början tyckte hon inte om hästen .
I början tyckte han inte om hästen .
Mina föräldrar tillät inte att jag gick ut med killar .
Den här maten var ju inte alls särskilt tokig !
På tv : n talar någon med allvarlig min om vårt lands framtidsproblem .
Ingen av dem deltog på mötet .
De använder teleskop för att betrakta himlen .
Jag hängde tavlan på väggen .
Vad skrattar du åt ?
Det säger sig självt att husdjur inte är tillåtna .
Skulle du kunna vara snäll och plocka ur diskmaskinen åt mig ?
Inga av de inbjudna gästerna har meddelat om de kan komma eller inte .
Vi kan kanske luncha någon annan dag .
Jag har bara femtio med rep .
Nu är det bra , varken för tungt eller för lätt .
Han köpte nya handskar .
Han iakttar varje liten rörelse jag gör .
Han stal pengarna i mitt kassaskåp .
Kan jag ta bilder här ?
Kan jag ta en bild här ?
Jag har en fråga .
Jag mutade polisen .
Tom och Mary paddlade kanot längs med floden sist jag såg dem .
Jag har alla de vänner som jag behöver .
De äter lunch i parken .
Jag är ingen häxa .
Är det där Tom ?
Skeppet syns fortfarande .
Båten syns fortfarande .
Du är den enda som jag kan lita på .
Han hade tre söner som blev advokater .
Jag värdesätter din vänskap högt .
Du är den ende som jag kan lita på .
Jag såg en vit hund hoppa över staketet .
Vem väntar du på ?
Han gav sin karriär som poet ett brått slut .
Datorn söker efter uppdateringar .
Tiden går för fort !
Jag blandar majonnäs med ketchup .
Man kan göra allt med majonnäs förutom att sitta på den .
Slottet var förfallet .
Hälsan är det viktigaste i livet .
En infraröd stråle består av elektromagnetisk strålning .
Jag vill ha två korv med bröd med mycket peppar .
Fattigdom lär en att äta bröd utan smör .
Tom tar en snabb joggingtur runt kvarteret varje morgon innan frukost .
Vad ska du göra under sommarlovet ?
Vad ska du göra på sommarlovet ?
Affären är öppen året runt .
Affären är öppen året om .
Jag ska inte göra illa dig .
Jag ska inte göra dig illa .
Jag är ingen nazist .
Hon översatte det ord för ord .
Hur svårt ska det vara egentligen ?
Han hade ingen anledning att gnälla på henne på det där sättet .
Mjölken kokade över .
Min mamma och jag är fullständigt olika .
Jag önskar att jag hade varit med henne då .
De kysste varandra .
Är du ledsen ?
Har du det bra ?
Vad ska du göra på fredag ?
Jag värdesätter vår vänskap .
Jag har inga nära vänner .
Jag är vacker .
Hunden rullade ihop sig i bädden .
Om jag bara kan stå på benen .
Det kan du inte säga .
De utgör att skickligt lag .
Ditt problem liknar mitt .
Jag kan inte rädda dig .
Jag var på bio .
Du måste vänta på nästa buss .
Jorgen älskar sin fru .
Norge heter " Norge " på norska .
Sverige heter " Sverige " på svenska .
Har ingen lärt dig att du inte får skolka ?
På högstadiet skolkade han dagarna i ända .
En person som skolkar kallas för skolkare .
Man kan inte bara skolka från skolan , utan från arbetet också .
Ett dussin ägg är färre än ett tjog .
När mörkret faller kryper tomtar och troll ut ur sina hålor i skogen .
Jag kan inte komma på texten .
De säger att han föddes i Tyskland .
Det sägs att han föddes i Tyskland .
Han har en Toyota .
Häng upp din kappa , tack .
Radion dog .
Han fjällade en fisk .
Han lämnade festen med bultande hjärta .
Jag måste få känna stadens puls .
Han försökte att inte vara allt för partisk .
Hon kunde inte låta bli att vara partisk i ärendet .
Orkanen skadade det lilla huset .
För henne är det en förolämpning .
Barnen knuffades .
Hon skickade ett brev till mig .
Hon skickade mig ett brev .
Har du någonsin sett en val ?
Du har två böcker .
Det kändes som om mitt ansikte brann .
Hon använder sällan nagellack .
Hennes nagellack hade börjat lossna .
Nia inte mig !
Finns det några biografer här i närheten ?
Jag tvättade bilen .
Ett äpple om dagen håller doktorn borta .
Hon satte sig på träningscykeln och trampade på tills hon blivit alldeles genomsvettig .
Jag behöver en anteckningsbok för att föra mina anteckningar .
Vad är skillnaden mellan amerikansk och brittisk engelska ?
Varför är ni alla här ?
Sent omsider gick det upp för mig att jag var ensam .
Ser du den mustaschprydda mannen där borta ?
Kan Tatoeba bidra till att rädda utrotningshotade språk ?
Engelska talas i många länder runt om i världen .
Hans mage skriker .
Hennes mage skriker .
Det är för kallt .
Den är för kall .
De stödde honom och hans politik fortfarande .
Han behöll hatten på .
Det är omöjligt att leva utan vatten .
Du är gammal nog att förstå .
Du är tillräckligt gammal för att förstå .
När kom Susana tillbaka ?
Vår lärare skrattar sällan .
Bob tittade förbi hos sin farbror .
Bilen förbrukar mycket bränsle .
Jag kunde inte ta mig utanför stadion på grund av folkmassan .
Ta väl hand om Tom .
Jag kan inte läsa franska , och ännu mindre tala det .
Jag funderar på att åka till Paris .
Jag kan inte förstå att jag precis sköt mig själv .
Tom kan tala flytande franska .
Tom kan tala franska flytande .
Tom kan prata flytande franska .
Tom kan prata franska flytande .
Vart gick pappa ?
Jag vill köpa en tjeckisk tröja .
Jag gjorde ett försök att simma över floden .
Vissa gillar kaffe och andra gillar te .
Vissa tycker om kaffe och andra tycker om te .
Vissa människor gillar kaffe och andra människor gillar te .
Vill du ha lite öl ?
Tack för alla dina kommentarer !
Han var siste man att komma fram .
Den här tanden sitter löst .
Jag kommer börja gråta !
Jag kommer börja grina !
Jane låtsades alltid att hon var väldigt rik .
Vill du ha någonting att äta ?
Vill du ha något att äta ?
Vill du ha nåt att äta ?
Jag gillar inte kvinnor utan personalitet .
Skådespelerskan har ett väldigt vackert namn .
Någon förstörde min kamera .
Någon gjorde sönder min kamera .
Någon hade sönder min kamera .
Jag skulle vilja ställa dig några till frågor .
Många träd tappar sina löv på vintern .
Många träd tappar löven på vintern .
Visade hon dig bilden ?
Visade han dig bilden ?
Vår engelsklärare lägger vikt vid uttalet .
Är inte det planen ?
Är det inte det som är planen ?
Han har skaffat sig vanan att stoppa händerna i fickorna .
Jag går till biblioteket två till tre gånger om veckan .
Jag går till biblioteket två eller tre gånger i veckan .
Jag går till biblioteket två till tre gånger per vecka .
Arbetsnarkomaner ser semesterdagar som slöseri med tid .
Arbetsnarkomaner ser semester som tidsslöseri .
Jag odlade tomater förra året och de smakade väldigt gott .
Jag odlade tomater förra året och de var väldigt goda .
Jag kan inte ta hennes plats som engelsklärare .
Ät dina grönsaker .
Han är en man att räkna med .
Han är en man som man kan räkna med .
Han sa åt eleverna att vara tysta .
Alla eleverna kommer från USA .
Han reste under antaget namn .
Han reste under fingerat namn .
Han reste under täcknamn .
Du måste återbetala dina skulder .
Ni måste återbetala era skulder .
Jag har skrivit ned alla siffror upp till trettioett .
Det är väldigt svårt att säga vilket land en person kommer ifrån .
Jag är på ett gräsligt humör i dag för jag har inte tillräckligt med pengar .
Jag fick reda på det av en ren händelse .
Bli inte sårad .
Tom är så där med alla .
Bli inte stött .
Tom är så där med alla .
De här skorna är gjorda i Italien .
Dessa skor är tillverkade i Italien .
Vi välkomnar alla som vill komma till festen .
Helens ord fyllde mig plötsligt med ny energi .
Helens ord fyllde mig plötsligt med ny kraft .
Hon är online flera timmar varje dag .
Jag var väldigt trött , så jag gick och la mig tidigt .
Du kan lika gärna säga det till honom i förväg .
Ni kan lika gärna säga det till honom i förväg .
Du låter besviken .
Ni låter besvikna .
De låter besvikna .
Det var lätt att hitta hans kontor .
Hon talar inte japanska hemma .
Hon pratar inte japanska hemma .
Han klär sig som en gentleman , men han talar och uppför sig som en clown .
Den här ölen är inte tillräckligt kall .
Den här ölen är inte kall nog .
I Europa och Amerika ser de hunden som en familjemedlem .
Ingen har lagt ned så mycket tid och ork i projektet som hon .
Det är ju inte direkt första gången som du kommer försent .
Den snälla systern hade bäddat in bäddsoffan lagom till att han kom fram .
Din otacksamhet är motbjudande .
Tom kan inte stå still .
Jag klarar inte av att se blod .
Jag klarar inte av synen av blod .
Jag står inte ut med tanken på att förlora Tom som vän .
Jag står inte ut med tanken på att förlora dig för evigt .
Jag klarar inte av sådana här filmer .
Jag klarar inte av sådan här musik .
Tom kan inte sjunga höga A.
Tom kan inte sjunga ett högt A.
Han har inte på sig en hatt .
Han har inte på sig hatt .
Han har inte hatt på sig .
Han har inte en hatt på sig .
Det är ett väldigt farligt system .
Nu är det dags för mig att krypa till kojs .
Jag tänkte krypa till kojs nu .
Jag önskar att vi hade mer tid .
Esperanto är talat i 120 länder runt om i världen .
Jag minns huset som jag växte upp i .
Öppna munnen .
Flickan har solglasögon .
Hon har solglasögon .
Han har solglasögon .
Efter filmen somnade de .
Mötet slutade klockan fem .
Skulle du kunna ögna igenom de där papperna lite ?
Min pappa kallar ibland stuprännor för " himlavattenavlägsningsrör " .
Min pappa röker .
Min far röker .
Jag skulle vilja att han vore här .
Problemet är inte så svårt att de skulle vara olösligt .
Jag vill ha tårta .
Jag måste påminna dig om ditt löfte .
Jag har samma problem som du hade .
Han var väldigt tålmodig .
Han hade ett väldigt tålamod .
Jag är ung .
Jag har ont i huvudet .
De dricker cola .
Han levde ett enkelt liv .
I år vill jag fira min födelsedag tillsammans med familj och vänner i Hagaparken .
De sökte alla efter det försvunna barnet .
De sökte alla det försvunna barnet .
Prata inte om det där framför honom .
Prata inte om det där i hans närvaro .
Prata inte om det där i hennes närvaro .
Öppna inte fönstret .
Jag skulle gärna tala med Judy .
De är inte alltid där .
Faktum är att hon läste inte ens brevet .
Dr .
Georges sekreterare är japanska .
Tom känner inte för att prata just nu .
De kämpade för religionsfrihet .
Jag förlorade allt .
Måndag börjar på söndag .
Jag studerade en stund i morse .
Jag pluggade en stund i morse .
Herr Smith har gjort det till en regel att ta en promenad varje morgon .
Vi kunde inte gå ut på grund av tyfonen .
Jag har precis varit på stationen för att vinka av min farbror .
Jag har precis varit på stationen för att vinka av min morbror .
Jag kysste henne på pannan .
Tom kysste Mary på pannan .
Hon kysste honom på pannan .
Han kysste mig på pannan .
Han kysste sin dotter på pannan .
Jag har sett en artikel på Tatoebabloggen om en ny version som ska komma ut snart .
Har du läst den ?
Hon gillar varken ormar eller matematik .
Hur är det med din syster ?
Det har varit ett dödsfall i din familj .
När jag hade packat färdigt min väska fick jag knappt igen den .
Du har tagit på dig hatten bakochfram .
De blev helt genomblöta i skyfallet .
Mary hjälpte sin mor att laga mat .
Mary hjälpte sin mamma att laga mat .
Tänk på vad du säger !
Lagom , tack !
Lagom är bäst .
Det enda svensken inte kan göra lagom är att fika .
Hon kommer hem igen lagom till jul .
Du tycker inte om mig .
Jag tycker om att lyssna på musik , speciellt jazz .
Har du tid att komma imorgon ?
Han kommer om en stund .
Var god och tag plats !
Ge mig en sked .
Ge mig skeden .
Jag väntar på dig på mitt rum .
Vad är Finlands huvudstad ?
Vilken är Finlands huvudstad ?
Tom fick Mary att gråta .
Söndag följs av Måndag .
Tom har inte hatt på sig varje dag .
Tom har på sig hatt varje dag .
Tom har på sig hatt nästan varje dag .
Tom har vanligtvis inte på sig hatt .
Tom har inte ofta på sig hatt .
Tom bär inte ofta hatt .
Tom har inte alltid hatt på sig .
Tom bär inte alltid hatt .
Tom har nästan aldrig på sig hatt .
Tom bär nästan aldrig hatt .
Tom har sällan på sig hatt .
Tom bär sällan hatt .
Sluta skjuta !
Vänta .
Skjut inte än .
Är det här Paris eller Marseille ?
Vill du ha lite äggröra ?
Du missbrukar dina maktbefogenheter .
Skulle du vilja ha lite äggröra ?
Tom äter ofta äggröra till frukost .
Din hund är där .
Din hund är här .
Er hund är här .
Lösenordet är " Muiriel " .
Jag tjänar 100 euro om dagen .
Jag saknar dig .
Det här är hans bil , tror jag .
Detta är hans bil , tror jag .
Ja , sa hon , du har rätt .
Hon är alltid kvick och slagfärdig .
Tom skrattar .
Tom har hemlängtan .
De vädrar alltid sängkläderna på torsdagar .
De bäddar ur sängen var tredje vecka .
De byter sängkläder var tredje vecka .
Tom är ostadig på benen .
Tom är vid sans .
En hunds nos är väldigt känslig .
Ett enormt monster är på väg ned från berget .
En man som inte spenderar tid med sin familj kan inte vara en riktig man .
En ponny är en liten häst .
En tredjedel är mindre än en halva .
Anpassning är nyckeln till överlevnad .
Sedermera antog han en ny identitet .
Jag gillar ris mer än bröd .
De hade inga skägg , inget hår och inga ögonbryn .
Vad kostar en öl ?
Snälla rätta mig när jag gör fel .
Alle man , överge skeppet !
Hela besättningen , överge skeppet !
En katt har en svans och fyra ben .
Ett DNA-test visade att han var oskyldig .
Tom håller på att kvävas .
Tom är vaken .
Tom blöder .
Tom är ensam .
Tom är uppmärksam .
Tom är alert .
Tom är bekymrad .
Tom är ängslig .
Tom är orolig .
Han skriver böcker .
Tom såg sig inte om .
Han är bög .
Jag tog ut kakan ur ugnen .
Världens snyggaste sambo fyller 25 i dag .
Han gillar indisk mat .
Aldrig prata med främlingar .
Hon är en långväga gäst .
Han tjänar tre gånger så mycket pengar som jag .
Han är tre år äldre än hon .
Hon är frånvarande för att hon är sjuk .
Födelsedagen firades med pompa och ståt .
Dimman lättnade .
Tack för att du accepterade min vänförfrågan på Facebook .
Vilken stor hund !
Och det här är min sida .
Och detta är min sida .
Hur länge har han varit borta ?
Hur länge har han varit frånvarande ?
Naturen är full av mysterium .
Min far tycker om starkt kaffe .
Sommaren är över .
I morgon ska jag gå och shoppa .
För länge sedan fanns här en bro .
För länge sedan fanns det en bro här .
Träffar du honom ofta ?
Träffar du henne ofta ?
Jag fick ta en veckas semester .
Jag har alltid en flaska mineralvatten med mig .
Han kom från Kanada för att träffa mig .
Hon kom från Kanada för att träffa mig .
Om du vill ha fred , förbered dig för krig .
George är väldigt pratsam .
Du har ett samtal .
Frukosten är färdig .
Jag har en hund som kan springa snabbt .
Detta barnet har växt upp normalt .
Jag tror inte att ungen kom till Tokyo själv .
Det är okej med mig .
Har du dina biljetter ?
Jag hoppas att något bra händer innan dagen är över .
Detta är väldigt lätt .
Min hund bet Tom .
Jag matade hunden .
Läs inte vad som är i brevet .
Bara ge det till Tom .
Jag tror han är ärlig .
Jag tror hon är ärlig .
Jag tror att hon är ärlig
Jag vet precis vem Tom tänker gifta sig med .
Folk ändras .
Det finns inte mycket du kan göra åt det .
Vem kommer att vinna i Ohio ?
Vem röstade du på ?
Vem blir den nästa presidenten av USA ?
Röstade du ?
John tände en tändsticka .
Du glömde att dividera med X här .
Vad gjorde han efter det ?
Vänta en sekund .
Detta telefonsamtalet kan vara viktigt .
Jag ska lära ut Esperanto i mitt land .
Jag är förföljd .
Dimman var så tjock att jag inte kunde se vart jag var påväg .
Ärligt talat , jag är inte särskilt imponerad av hans idée .
Jag svär att jag aldrig ska göra det igen .
Är han inte söt när han är arg ?
Jag skrattade väldigt mycket när jag såg det där .
Tom brukade röka två paket cigaretter varje dag .
Tom spenderade hela dagen med att designa en hemsida åt en ny kund .
Har du blivit en ängel ?
Vill du ha te eller något ?
Jag sovde väldigt bra .
Mitt te är för sött .
Vi hade rätt .
Hur träffade du din partner ?
Jag tvättade min T-shirt .
Släpp ankaret !
Ju mer pengar vi har , desto mer vill vi ha .
Hur var din dag idag ?
Hon är så jävla charmig !
Visa hur man gör det där .
Visa mig .
Tom alltid på sig en hatt .
Tom har nästan alltid på sig en hatt .
Tom har ofta på sig en hatt .
Tom har ibland på sig en hatt .
Jag glömde min egen födelsedag .
Faktiskt så hittade jag på det där .
Faktiskt så är jag inte särskilt säker .
Kan du tro att detta faktiskt händer ?
Hände det verkligen ?
Sa verkligen Tom det ?
Trodde du verkligen det ?
Läste du verkligen det ?
Gav du verkligen Tom pengar ?
Såg du verkligen Tom ?
Jag jobbar faktiskt här .
Jag gick faktiskt aldrig på högskola .
Jag såg det faktiskt inte själv .
Jag trodde inte att Tom faktiskt skulle prova det .
Jag har faktiskt aldrig träffat Tom .
Jag såg det faktiskt aldrig .
Jag är faktiskt en väldigt bra förare .
Jag är faktiskt ganska seriös .
Jag har faktiskt kul ikväll .
Jag är faktiskt ganska trött .
Jag är faktiskt väldigt lycklig .
Jag är faktiskt här för att hjälpa dig .
Jag har faktiskt aldrig varit full .
Jag är faktiskt väldigt upptagen .
Jag har faktiskt aldrig spelat golf .
Händer detta verkligen ?
Det är faktiskt inte riktigt så enkelt .
Det var faktiskt inte så illa .
Det låter som om du faktiskt menar det .
Det var faktiskt mitt fel .
Det är faktiskt mycket enklare än vad det ser ut .
Det är faktiskt en bra poäng .
Det är faktiskt inte sant .
Det är faktiskt ganska smart .
Det är faktiskt bra nyheter .
Det är därför jag är här , faktiskt .
Tom trodde faktiskt på dig .
Tom gjorde faktiskt det han sa att han skulle göra .
Detta är total demagogi .
Alla dörrar i huset var stängda .
Tom kom faktiskt på det själv .
Tom fick faktiskt Mary till att dansa med honom .
Tom gillar faktiskt Mary .
Tom spelar faktiskt inte mycket .
Tom pratar faktiskt inte mycket Franska .
Tom är faktiskt väldigt bra på att laga mat .
Tom var faktiskt inte där .
Toms party var ganska roligt , faktiskt .
Jag har inga kläder att använda .
Jag har inga rena kläder att använda .
Snälla gå ut härifrån genast .
Snälla gå ut ur mitt kontor genast .
Jag kan inte låta dem fånga mig .
Jag kan inte låta dem fånga dig .
Vem var det som faktiskt genomförde operationen ?
Vi behöver faktiskt inte göra det nu .
Jag har ingenting att läsa .
Jag har inga böcker att läsa .
Jag har inget att skriva med .
Jag har ingenstans att gå .
Jag behöver förstå vad denna mening betyder .
Vi gick ut på en promenad efter frukost .
Han är inte alltid glad .
Öppna inte lådan än .
Öppna inte presenten än .
Varför svarar du inte ?
Jag tror inte att kärlek finns .
Jag kan inte ens göra en omelett .
Jag kan inte förstå någonting av det han säger .
Han gick upp tidigt för att han skulle komma i tid till tåget .
Du ska alltid skydda dina ögon från direkt solljus .
Att bli klar med detta jobbet innan tisdag kommer att vara enkelt .
Han gillar grönsaker , framförallt vitkål .
Det vore bättre om du inte åt innan du gick till sängs .
Kan du snälla säga hur lång du är och din vikt ?
Kan du snälla säga hur lång du är och hur mycket du väger ?
Snälla ge mig ett plåster och lite medicin .
Jag mår inte bra .
Snälla ge mig lite medicin .
Min far har slutat röka på grund av sin hälsa .
Min far har slutat röka för sin hälsas skull .
Tom sa alltid att han ville lära sig spela mahjong .
Toms mamma sa alltid till honom att han borde äta mer grönsaker .
Du kanske har rätt .
Det var väldigt roligt .
Det var riktigt roligt .
Det var hemskt roligt .
Det var extremt roligt .
Det var ganska roligt .
Det var nästan roligt .
Det var inte roligt alls .
Klockan är nästan sju .
Vi måste gå till skolan .
Jag har fyra datorer , men två av dem är så gamla att jag inte använder dem längre .
Toms fru gillar inte när han röker i vardagsrummet .
Jag är riktigt trött .
Idag gick jag alldeles för mycket .
Ljudet väckte mig från min sömn .
Ljudet kommer att väcka bebisen .
Ingen kunde förklara hur saken var gjord .
Fången var bakom galler i två månader .
Satte du på frimärket på brevet ?
Varför provade du inte klänningen innan du köpte den ?
Rummet är fullt av folk .
Min bror och jag delade rummet .
Jag hittade rummet tomt .
Har rummet ett badkar ?
Rummet städas av fru Smith .
Rummet kommer att målas imorgon .
Det var en massa möbler i rummet .
Det fanns ingen i rummet .
Rummet har två fönster .
Det fanns nästan ingenting i rummet .
Det finns ett piano i rummet .
Det finns en TV i rummet .
Det finns två hundra personer i rummet .
Damen förblev tyst .
Damen är över åttio .
Paret hade ett lyckligt liv .
Fyll flaskan med vatten .
Den stackars mannen blev äntligen en känd artist .
Den sjuka mannens liv är i fara .
Sjukhuset öppnade förra månaden .
Isen är väldigt tjock .
Ord kan inte beskriva skönheten .
Den vackra kvinna är vänlig .
Planet flög över Mt .
Fuji .
Planet gjorde en perfekt landning .
Det var femtio passagerare på planet .
Dörren öppnar nu .
Dörren är öppen nu .
Tjejen är ensam .
Jag är säker på att jag rätt nummer .
Det var väldigt kallt den kvällen .
Jag kan inte stå ut med ljudet .
Ta bort lådan .
Titta inte in i lådan .
Lådan är för tung för att lyftas .
Lådan är nästan tom.
Lådan var nästan full .
Det är en massa ägg i lådan .
Lägg ingenting på lådan .
Vad finns i lådan ?
Det fanns ingenting i lådan .
Lådan var full av böcker .
Du måste lära dig engelska , vare sig du vill det eller ej .
Du måste lära dig engelska , vare sig du vill det eller inte .
Han blev blind .
Han blödde näsblod .
Klä på dig .
Vänta inte .
Stanna inte .
Stirra inte .
Sjung inte .
Spring inte !
Rör dig inte !
Han klarade det .
Han gick hem .
Han promenerade hem .
Han ser stark ut .
Tom är trött .
Tom är konstig .
Tom är hög .
Snälla lämna .
Du ser precis ut som din pappa .
Han har aldrig varit i Amerika .
Jag har inte tid att läsa böcker .
Jag behöver mer tid .
Kan du japanska ?
Jag kommer att behöva din hjälp .
Jag vill inte prata om det .
Han vill inte prata om det .
Hon pratade aldrig om det .
Han pratade aldrig om det .
Hon är ganska söt .
Vad för fråga är det där ?
Gillar du sött te ?
Skulle du ha något emot att jag ställer en fråga ?
Du frågar ofta frågor som jag inte kan svara på .
Snälla fråga inte en sådan fråga .
Låt mig fråga en fråga .
Jag ville bara ställa en fråga .
Jag ställde inga frågor .
Fråga inte , bara gör det .
Har du lärt dig din läxa ?
Det är hemligt .
Vad vill du ?
Vem åt den sista kakan ?
Ställ inga frågor .
Vad gjorde du i skolan idag ?
Ingen står över lagen .
Tom är elak .
Tom är fet .
Tom är döv .
Tom är uttråkad .
Tom har fel .
Är den vit ?
Jag behöver er .
Han springer .
Han sprang .
Gå iväg .
Jag också .
Tvätta dig .
Ha det så roligt .
Jag förstår .
Jag använder det .
Får jag öppna en burk ?
Mina ögon är ömma .
Min far är inte hemma .
Min näsa kliar .
Gör ditt val .
Vad gjorde Jean ?
Vad har hon ?
Vad är det Ken äter ?
Vad är det där borta ?
När börjar det ?
Var gör det ont ?
Jag gillar den personen .
Var är ditt rum ?
Vart ska vi gå ?
Tom kände sig väldigt ensam .
Tom har en liten paj .
Tom har många talanger .
Tom är en bra person
Tom kommer aldrig i tid .
Tom slog ner honom .
Tom ser väldigt glad ut .
Håll dig undan från hunden .
Gå inte nära hunden .
Ligg på din högra sida .
Marias hår är långt .
Mary gillar att titta på TV .
Kan jag ställa ner den här ?
Morfar köpte den till mig .
Har du ätit lunch än ?
Har du någonsin varit på TV ?
Har du matat hunden än ?
Ge mig en flaska vin .
Mary och Jane är kusiner .
Mary gillar mjölk väldigt mycket .
Min lägenhet är i närheten .
Min far älskar min mor .
Min far är duktig på att simma .
Min katt dog igår .
Var är Toms klassrum ?
Vart skulle du vilja åka ?
Min far är stolt över det faktum att han aldrig varit i en trafikolycka .
Vem vill du prata med ?
Vem är det som äger pistolen ?
Vem mer kom till festen ?
Varför är du arg på honom ?
Varför ser du så ledsen ut ?
Varför är du så trött idag ?
Varför gjorde han en sån sak ?
Mary sprang .
Stå upp .
Ursäkta mig .
Jag kan springa .
Jag kan åka skidor .
Jag ger upp .
Släpp in mig .
Självklart !
Självklart .
Det är okej .
Försök igen .
Vem vet ?
Har jag fel ?
Mår du bra ?
Fåglar sjunger .
Får jag hjälpa ?
Han är snäll .
Jag kan simma .
Jag gillar honom .
Jag älskar henne .
Jag betalar .
Jag är upptagen .
Jag är ledig .
Är det gratis ?
Släpp ut mig !
Låt mig betala .
Låt mig se .
Titta på mig .
Ta en buss .
Prata med mig !
Vi är män .
Du kan gå .
Gråt inte .
Han får komma .
Han ljuger .
Hur mår Mary ?
Jag är längre .
Jag gillar båda .
Jag gillar jazz .
Jag älskar rock .
Jag försov mig .
Jag blev avskedad .
Jag var trött .
Jag är vaken .
Jag är pank .
Jag har rätt .
Min lägenhet ligger här i närheten .
Förlåt .
Livet är roligt .
Snälla kom .
Jag är mänsklig .
Jag är människa .
Jag är en människa .
Hur uttalar man ditt namn ?
Hur uttalas ditt namn ?
Mina bröder skämtar alltid .
Ingen av hans elever kunde lösa uppgiften .
Ingen av hennes elever kunde lösa uppgiften .
Alla skrattade åt hans misstag .
Alla skrattade åt hennes misstag .
Han har säkert rätt .
Hon har säkert rätt .
Katten satt på bordet .
Att blir klar med det här jobbet innan tisdag kommer att bli enkelt .
Att bli klar med det här jobbet innan tisdag kommer att vara enkelt .
Att bli klar med detta jobb innan tisdag kommer att bli enkelt .
Att bli klar med detta jobb innan tisdag kommer att vara enkelt .
Kaffe eller te ?
Jag tycker att esperanto är mycket svårt .
Stationen ligger nära hotellet .
Vet du varför himlen är blå ?
Det där gjorde du med flit !
Följ efter den där bilen .
Mamma vaknar genast när man kittlar henne under fötterna .
Hon bet honom .
Hon slog honom .
Hon är snäll .
Gillar du den här trädgården ?
Gillar du denna trädgård ?
Tycker du om den här trädgården ?
Stäng av den .
Tycker du om denna trädgård ?
Hade jag fel ?
Tom hyser stor respekt för Mary .
Hur är läget ?
Vad händer ?
Alice log .
Är du vilse ?
Kan du komma ?
Kom med oss .
Prata inte !
Han har en bil .
Han älskar henne .
Han var själv .
Han var ensam .
Han var modig .
Han är smart .
Han är intelligent .
Jag åt kaviar .
Jag har en penna .
Jag gillade Tony .
Jag kommer .
Är det sant ?
Det var natt .
Det är min CD-skiva .
Det är min CD .
Mary kom in .
Ingen vet .
Snälla ta det lugnt .
Snälla lugna ner dig .
Hon är lycklig .
Hon är tystlåten .
Hon är tyst .
Hon känner mig .
Hon gick ut .
Det är mitt .
Den är min .
Du är sen .
Du är inte i tid .
Han kramade henne .
Han är stark .
Tom skynda dig .
Jag tror på dig .
Jag gillar vinter .
Jag såg ett flygplan .
Jag sålde en bok .
Jag använder Firefox .
Jag var hemma .
Jag är säker .
Jag är hälsosam .
Jag är seriös .
Jag är så mätt .
Jag är utsvulten .
Det är molnigt .
Det är måndag .
Det är mitt jobb .
Hör av dig !
Mary kan simma .
Får jag gå hem ?
Hon undviker mig .
Hon kom sist .
Hon blev arg .
Hon hatade honom .
Hon hatar honom .
Hon hjälper honom .
Hon gråter .
Hon gillar honom .
Hon ser ledsen ut .
Hon älskar honom .
Hon älskar Tom .
Hon var modig .
Hon gick hem .
Tom är frånvarande .
Vad är detta ?
Var är du ?
Kommer hon att komma ?
Du ser upptagen ut .
Du ser sjuk ut .
Du borde gå .
Var inte ledsen .
Varför är tjejer så komplicerade ?
Tjejer är inte komplicerade .
Män är simpla .
Du lovade ju att komma hem till sommaren .
Jag har ingen CD-spelare men jag köpte CD-skivan i alla fall .
Pengar är roten till allt ont .
Jag förstår inte vad det är han vill ha .
Jag ber så hemskt mycket om ursäkt , men jag jag måste be om att få ändra datumet för mötet till 6 mars på grund av personliga skäl .
Jag går alltid till skolan till fots .
Han oroar sig över testresultatet .
En del av äpplena som låg i lådan var ruttna .
Jag skäms över att jag sade det på det sättet .
Sam lovade att betala i slutet av månaden .
Jag sökte skydd från regnet under den affärens tak .
Hon hoppade på tunnelbanan i Ginza .
Min familj jobbar fortfarande så det dröjer fortfarande innan de kan åka till Texas .
Jag saknade min familj , så jag återvände hem .
Om jag har fått jobb till nästa år och kan ta ledigt i en längre period så åker jag snart till Japan !
Jag skulle uppskatta om ni kunde komma .
Det här stället är inte så nytt , men på plussidan så kan man grilla på verandan och hyra en portabel stekplatta för 2000 yen .
Är det OK om vi inte åker till Costco den här gången ?
Planen är att jag ska ha slutat mitt jobb då , så jag kanske kan gå !
Jag var säker på att du skulle stanna i Japan längre än så .
Jag kommer inte vara hemma från morgonen så jag kan inte kolla min mejl på PC : n så skicka till min mobil istället .
Aichis stränder är inte särskilt vackra .
Det blir lite svårt för mig att åka till Europa , men om ni har någon tillställning i Japan så vill jag gärna gå !
För mig så blir det för första gången på ett bra tag som jag inte åker hem till Hokkaido för att fira nyår .
Det finns bara två primtal mellan 10 och 14 .
Det är många som faktiskt är för att införa dödsstraff .
Det är uppenbart att korruptionen är ett stort problem .
Det ser ut att bli ett lovande år för det svenska modeundret .
Själv föredrar jag vodka , men jag har inget emot att ta en likör ibland .
Jag tillbringade en helg i New York , men gosse vad jag hatade det .
Det blir till att köpa en ny vinterjacka snart .
Jag insåg just att jag har haft den här i snart 6 år .
Min flickvän är helt tokig i Forever 21 , men det är åtminstone billigt .
Det är helt löjligt hur mycket pengar vissa sitter på .
Skit också , jag glömde att ställa tillbaka smöret i kylskåpet .. !
Jag förstår inte vad det är med den här osten , den började lukta skunk bara efter en vecka .
Man var tvungen att först stå i kö för att få en en lapp där det stod när man skulle få ställa sig i den riktiga kön .
Jag har aldrig varit med om något liknande .
Japans varma källor kan visa sig vara en viktig energikälla .
Min fru slår mig .
Varje gång jag sätter på mikrovågsugnen så slutar mitt Wi-Fi att fungera , det är extremt irriterande .
De kommer bli de första som ställs mot väggen när revolutionen kommer .
Johannes tycker inte om när man använder begrepp som " ras " .
Hur många skyskrapor finns det egentligen i Shanghai ?
Robert anmälde sig till någon sliskig dokusåpa av något slag , men som tur var gick han inte vidare .
Från mitt fönster har jag en kvintessentiellt japansk utsikt .
En god mandellikör skulle allt sitta bra nu .
Nej , jag har väl inte sagt att jag har något emot homosexuella heller ?
Det är uppenbart att moderaterna inte står högt i kurs bland studenterna på Smålands nation .
Jag skulle vilja säga att det är så att det är stockholmare som har svårt med folk från landsbygden , snarare än tvärtom .
Det är nog inte många som föredrar Uppsala framför Lund .
Det tog bara några veckor innan utbytesttudenterna råkade i luven på varandra .
Hellre död än röd .
Hjärtat sitter till vänster .
Mobbning är så klart ett allvarligt problem , men samtidigt måste vi inse att en nollvision här är omöjlig .
Många tyckte att Arne var lite för intim med sina elever .
Det fanns till och med dem som sa att han " kladdade " .
Det förekommer så mycket rasistiska kommentarer i svenska tidningars kommentarsfält att jag inte längre ids bry mig .
Jag har inte bett om någon jävla hjälp , det ska du ha klart för dig !
Det ska du ha jävligt klart för dig !
Visst , min mamma är prostituerad , men på den ljusa sidan så har vi åtminstone någonstans att bo .
Det skulle aldrig ens falla mig in att påstå något sådant .
Robotarna kommer att ta över en dag , det kan du vara säker på .
Usch , vilket klantarsel din far är .
Men skit på dig då , din jävla idiot .
Visst älskar jag Finland , men jag står inte ut med finnarna .
Du kanske inte tittar så mycket på TV ?
Man får nog leta både länge och noga om man överhuvudtaget ska ha en chans att hitta en mer klentrogen man än din farbror .
Din mamma är en riktig snuskhummer , Pelle .
Jag orkar inte med hennes insinuationer !
Det är väl inte svårare än att klart och tydligt säga " nej " .
Hon har inte mycket till skrupler , din mormor .
Bra jobbat , gubbar .
Det finns nog inte många som överhuvudtaget har något positivt att säga om SJ .
Om jag fick bestämma skulle man släppa en mindre atombomb över SJ : s huvudkontor i Stockholm och sen börja om på ny kula .
Om tåget inte är försenat än , så kommer det att bli det snart .
Tids nog ska nog även detta tåg bli försenat .
Jag har fått nog av alla dessa kissnödiga kvällstidningskrönikörer .
Håll ett öga på Tom .
Hon såg mer vacker ut än någonsin förrut .
Kan jag räkna med dig ?
Kan jag lita på dig ?
Jag är riktigt stolt över dig .
Jag skulle vilja ha ett ord med dig .
Jag antar att vi har gjort ett helt okej jobb eftersom ingen har klagat .
Vill du att jag ska ringa polisen ?
Jag blev så ställd att jag började gråta .
Min man blev så ställd att han tappade sina bilnycklar .
Jag har inte mycket till övers för Hollywoods superhjältefilmer .
Varför återkommer Hollywood ständigt till dessa män i trikåer ?
Du kan kalla det för dialektalt bäst du vill , jag är övertygad om att det är ett rikssvenskt uttryck .
Min mamma är svensklärare så hon överreagerar så in i vassen så fort man råkar använda ett lite svengelskt uttryck .
Min far är faktiskt universitetslektor , så vet hut .
Jag vet att jag kan verka lite slemmig , men jag kan faktiskt vara ganska hårdför .
Det är nog mycket få som skulle få för sig att uttrycka sig på det sättet framför en statsminister .
Kommer du hit ofta ?
Det var väl bara det som fattades , nu har min dotter en bulle i ugnen också !
Fåntratt !
Man kan inte multiplicera så här stora tal för hands !
Ankdamma mig hit och ankdamma mig dit , jag tycker inte att det är något fel på debatten .
Men det var väl ett evinnerligt tjat !
Nej , du får ingen snickers !
Ja , så kan man väl tycka , om man nu vill .
Sicken retsticka , va !
Kom inte här och tro att du är något .
Visst kan du kalla mig för idiot .
Vad vill du jag ska säga , det är sån musik som jag gillar .
Jag håller inte med , det är inte rasistiskt att använda ordet " ras " .
Skynda på med inhalatorn , Jocke håller på att få ett astmaanfall !
Nej , nej och åter nej .
Oj , en sverigedemokrat uttryckte sig rasistiskt , stoppa pressarna !
Det finns ju vissa uttryck som numera bara används ironiskt .
Ingen har bett dig att hålla med , men du kan väl åtminstone acceptera att det finns personer som har andra åsikter än dig ?
Fet chans .
Jaha , det var ju just en stor överraskning också .
Nä , säger du det ?
Du , intresseklubben antecknar .
Men har du svårt att förstå eller låtsas du bara ?
Bara så du vet : det är ingen som tycker synd om dig .
Jag har en farbror som bor i Provence , han är helt lyrisk över bouillabaissen de har där .
Gå och häng dig , apjävel !
Visst kan det vara traumatiskt , men än sen ?
Jag litar inte på politiker .
Min pappa sade alltid att socialdemokrater har en smuts som inte går bort , i själen .
Min mamma brukade säga att det inte finns någon som har mindre medlidande än en moderat .
Båda mina föräldrar var arbetslösa , men det hindrade dem inte från att ta väl hand om mig och mina 23 syskon .
Snubben som står i hörnet där borta kan röka upp en cigarett på mindre än en minut .
På 80-talet var det minsann andra bullar som gällde .
Men det var väl mig ett jävla tjat om den förbannade 30-talsjazzen !
Jag tar en kebabpizza special , med blandad sås .
Jag tänker under inga omständigheter låta dig ta över min fars rederi .
Detta rederi ska då aldrig falla i en göteborgares händer !
Det brinner i rederiet !
Många grekiska skeppare förmodas lämna landet om en sådan reform förs igenom .
Jag trodde att jag gjort klart för dig att detta rederi inte är till salu !
Min far ville att min äldre bror skulle ta över rederiet , men tji fick han .
Det här är ett familjerederi och vi kommer aldrig att sälja det !
Trevligt varuhus , vore ju synd om något skulle hända det ...
Hur fan kan man få för sig att sitta och äta varmkorv på toaletten ?
Hur är din farsa funtad egentligen ? !
Man gör väl inte direkt sina läsare en tjänst genom att kalla detta parti för reformvänligt .
Svårt att tro , men så är det .
Förlåt mig , jag har bråttom , måste iväg nu illa bums !
Du såg hunden som tillhör den man som jag flirtade med .
Driver du med mig ?
Du måste skämta !
Ge det till henne .
Ge den till henne .
Ge den till honom .
Ge det till honom .
Har du ätit ?
Han är en författare .
Han ser ung ut .
Verkar som om han är trött .
Han var hemma .
Jag åt för mycket .
Jag ogillar ägg .
Jag bryr mig inte .
Jag har inget emot det .
Jag har en idé .
Han sprang så fort som han förmådde .
Vi ska på bio .
Kom med .
Vi hyrde lägenheten .
Han fäste affischen på anslagstavlan med häftstift .
Vad gjorde du i går kväll ?
Tom gjorde det , eller hur ?
Vad sägs om att sätta på en kopp te ?
Hon föreslog för honom att resa utomlands medan han fortfarande är ung .
Det var en incident förra året med en säkerhetsvakt som avlossade ett vådaskott inne på en toalett .
Jag är färdig .
Jag måste köpa en .
Jag reser ofta .
Jag såg henne simma .
Jag kommer inte att förlora .
Jag är en doktor .
Jag är upptagen nu .
Jag är så lycklig .
Jag är jättetjock .
Är han från Japan ?
Är hon hemma ?
Lämna mig ifred !
Låt mig vara !
Låt mig vara .
Lämna mig ifred .
Lyssna på detta !
Lyssna !
Lynn springer snabbt .
Många fiskar dog .
Mr .
Smith kom .
Säg det tydligt .
Sluta göra omsvep och kom till saken .
Sluta gå som katten kring en het gröt och kom till saken .
Vad saknas ?
" Vill du lämna ett meddelande ? "
" Nej , tack . "
" Han har varit sjuk . "
" Jaså , jag hoppas att det inte är någonting allvarligt . "
En man som kan två språk är värd två män .
En förbipasserande bil körde i en vattenpöl och stänkte ned hela mig .
En sexsiffrig inkomst är inte ovanligt för en läkare .
Tom är skyldig .
Hon kom ensam .
Hon lurade honom .
Hon hjälpte honom .
Hon kramade honom .
Hon är en sjuksköterska .
Hon är ute nu .
Hon sparkade honom .
Hon kysste honom .
Hon älskar katter .
Hon saknar honom .
Hon sjunger bra .
Han är bra på att sjunga .
Ta din tid .
Det stämmer !
Det är sant .
Korrekt !
Det är konstigt .
De hatade Tom .
De bråkade .
Detta är min bil .
Tom ser blek ut .
Tvätta ditt ansikte .
Var ligger Paris ?
Var är Tony ?
Vem förstörde denna ?
Vem förstörde det här ?
Varför frågar du ?
Varför ljuger du ?
Tråkar jag ut dig ?
Skämtar du ?
Skämta inte med mig !
Städa ditt rum .
Känner du henne ?
Känner du honom ?
Känner du igen honom ?
Vet du vem hon är ?
Ge inte upp !
Kör försiktigt .
Följ den bilen .
Har han kommit än ?
Ha en bra dag .
Han har gått ut .
Han har tio kossor .
Han har tio kor .
Han är ogift .
Han gillar att springa .
Hon gillar att springa .
Han blev av med sitt jobb .
Han älskar tåg .
Han studerar .
Han pluggar .
Snälla hjälp mig .
Hur är det med din pappa ?
Hur mår din pappa ?
Jag köpte en bok .
Jag hatar politik .
Jag avskyr politik .
Jag har två bilar .
Jag bor i Japan .
Jag behöver någon .
Han spelade tennis .
Jag brukade spela tennis .
Jag spelade tennis .
Jag springer varje dag .
Jag joggar varje dag .
Jag vill ha en gitarr .
Jag vill ha den väskan .
Jag vill sova .
Jag är nöjd .
Jag är belåten .
Jag är väldigt upptagen .
Jag kom på det .
Är någon hemma ?
Andas han ?
Är hon Japansk ?
Det kommer inte att funka .
Det kommer inte att gå .
Jag bjuder .
Det är för högt .
Den är för stor .
Den är väldigt stor .
Kate är förkyld .
Låt mig se det där .
Titta bakom dig .
Min hat trillade av .
Öppna flaskan .
Tatoebaprojektet , som återfinns online på tatoeba.org , går ut på att skapa en stor databas med exempelmeningar översatta till många språk .
Hörde du det där ?
Fråga Tom .
Ta det lugnt .
Var trevlig .
Kom igen .
Hämta Tom .
Sluta !
Lägg av !
Var still .
Stilla .
Kör vidare .
Ducka .
Fortsätt in .
Hugg tag i Tom .
Blidka mig .
Gör mig till viljes .
Låt det vara .
Låt den vara .
Lämna mig .
Lämna oss .
Gift dig med mig .
Använd den här .
Använd det här .
Använd denna .
Använd detta .
Varna Tom .
Se på mig .
Titta på oss .
Se på oss .
Skriv till mig .
Sikta .
Skjut !
Lugna dig .
Dö inte .
Ta tag i den där .
Flytta på dig .
Sluta med det där .
Sluta upp med det där .
Ryck upp dig .
Skynda dig !
Spring för livet !
Gör det inte .
Gå inte .
Han låtsas .
Låt mig hjälpa till .
Tom är död .
Ringde Tom ?
Har Tom ringt ?
Ser jag OK ut ?
Ser jag bra ut ?
Ta dig ett glas .
Ta en drink .
Han är så söt .
Hur går det med skolan ?
Hur går det på skolan ?
Hur går det i skolan ?
Jag måste gå .
Jag drog mig ur .
Jag klarar mig .
Jag kommer att vara här .
Jag är här .
Jag stannar här .
Jag fixar en .
Jag hämtar en .
Jag ska betala dig .
Jag fick dig .
Jag har dig .
Peka ut den .
Peka ut det .
Hon gillade det .
Hon gillade den .
Hon tyckte om det .
Hon tyckte om den .
Stanna bilen .
Tom hatar mig .
Tom behöver mig .
Tom ryckte på axlarna .
Vi kommer överens .
Vi kommer väl överens .
Du är konstig .
Gjorde jag det där ?
Var det jag som gjorde det där ?
Gör det snabbt .
Gör det fort .
Vet Tom ?
Vet Tom om det ?
Var inte elak .
Var inte oförskämd .
Var inte ohövlig .
Var inte ohyfsad .
Gör inte det här .
Gör inte detta .
Var inte uppkäftig .
Var inte kaxig .
Han är irriterande .
Han är besvärlig .
Hur illa är det ?
Jag kan inte dansa .
Jag gjorde ingenting .
Jag går först .
Jag kommer att gå först .
Jag kommer att hjälpa dig .
Jag ska berätta för dig .
Jag kommer att berätta för dig .
Jag berättar för dig .
Jag är bara lat .
Mary är konstig .
Ta det i din egen takt .
Hon är grym .
Ta bara en .
Det är en plan .
Det är mycket .
Det här är konstigt .
Detta är konstigt .
Detta är underligt .
Det här är underligt .
Tom hatar dig .
Tom är en sportig typ .
Tom är en idrottare .
Tom är en idrottskille .
Tom är inte rolig .
Tom är rädd .
Tom släppte in mig .
Tom hade rätt .
Var Tom ensam ?
Vi kan inte misslyckas .
Vi måste gå .
Vi borde äta .
Vi förstår .
Vi ska vi göra ?
Vad ska vi ta oss till ?
När var det ?
Du är en snobb .
Du är inte rolig .
Kommer jag att dö ?
Är vi vänner ?
Gråter du ?
Grinar du ?
Kan jag komma med dig ?
Kan jag sitta ned ?
Hallå , är det någon där ?
Herregud , vilken tid det tar !
Jo , visst kan jag göra det .
Han träffade sin älskling på restaurangen .
Tänk , vad fort tiden går .
Släpp tag i min arm !
Ser du killen där borta med svart jacka ?
Oroa dig inte över sådana småsaker .
En miss till och du är ute .
Tack , det räcker .
Tjena , grabben !
Håll dig bara lugn så kommer allt att gå bra .
Jaså , vem har sagt det ?
Jag ska träffa en kompis efter skolan .
Stick härifrån !
Nu sticker vi .
Välkommen till vår enkla boning .
Mina herrar och damer , låt mig presentera …
Kan du fixa den här åt mig ?
Skjut inte !
Kom tillbaka hit .
Fattade du ?
Provade du det ?
Känner vi dig ?
Känner vi er ?
Lovar du ?
Lovar ni ?
Spelar det någon roll ?
Bryr du dig inte ?
Sov lite .
Har du sovit ?
Han fick jobbet .
Bromsa .
Hur illa var det ?
Hur dåligt var det ?
Hur kan jag hjälpa till ?
Hur kan jag hjälpa ?
Hur var Hawaii ?
Jag ringde i förväg .
Jag kan hjälpa dig .
Jag gjorde det inte .
Jag hörde röster .
Jag träffade honom precis .
Jag behöver min jacka .
Jag behöver min rock .
Jag behöver min kappa .
Jag sa stick .
Jag tar den .
Jag ska göra det nu .
Jag ska ta hand om det .
Jag tar hand om det .
Jag betalar extra .
Jag ska betala extra .
Jag kommer att betala extra .
Jag ska skjuta dig .
Jag skjuter dig .
Jag kommer att skjuta dig .
Jag väntar här .
Jag kommer att vänta här .
Jag älskar ditt hår .
Jag tar aldrig sovmorgon .
Jag föredrar att gå .
Jag såg allt .
Jag tror att Tom gick .
Jag skulle vilja hjälpa till .
Jag kommer att vara hos Tom .
Jag är hos Tom .
Jag ska kolla igen .
Jag ska hämta min jacka .
Jag ska ta min jacka .
Jag ska hämta min rock .
Jag ska ta min rock .
Jag ska hämta min kappa .
Jag ska ta min kappa .
Jag hämtar mina nycklar .
Jag hämtar nycklarna .
Jag ska hämta mina nycklar .
Jag ska hämta nycklarna .
Jag hämtar bilen .
Jag ska hämta bilen .
Jag ska gå och handla .
Jag ska gå och shoppa .
Jag följer med dig .
Jag kommer att följa med dig .
Jag ska följa med dig .
Jag tar hand om det här .
Jag kommer att ta hand om det här .
Jag ska ta hand om det här .
Jag hämtar upp Tom .
Jag kommer att hämta upp Tom .
Jag ska hämta upp Tom .
Jag pratar med Tom .
Jag ska prata med Tom .
Jag kommer att prata med Tom .
Jag är redan rik .
Finns det något godare än kladdkaka och glass ?
Kladdkaka och glass kan vara det godaste som finns .
1,6 mil är inte en kort sträcka .
16 kilometer är inte en kort sträcka .
Jag ska försöka .
Jag kommer att försöka .
Jag är på vinden .
Jag är på vindsvåningen .
Jag är ingen tiggare .
Jag är trött på det här .
Jag har fått nog av det här .
Det är din rättighet .
Det fick mig att skratta .
Mary knäböjer .
Snälla kör in till trottoarkanten .
Så vad hände ?
Sluta plåga mig .
Sluta tjata på mig .
Ta hand om Tom .
Det är gammal skåpmat .
Bucklan var min .
Pottan var min .
Krukan var min .
Burken var min .
Kannan var min .
Grytan var min .
Haschet var mitt .
De kommer med undanflykter .
De slingrar sig .
De överstegrar .
De kör fast .
Det här är inte rätt .
Detta är inte rätt .
Detta stämmer inte .
Det här stämmer inte .
Tom frågade ut mig .
Tom åt sig mätt .
Tom åt så mycket han orkade .
Tom studsade tillbaka .
Jag är musiker .
Jag är arg på dig .
Jag är precis här .
Låt mig hämta Tom .
Visa oss runt .
De där är trevliga .
De där är fina .
Tom kan inte komma .
Tom kan inte stanna .
Tom kan inte gå .
Tom klappade ihop .
Tom tog knäcken på sig .
Tom dog ensam .
Tom är ett äckel .
Tom är en hippie .
Tom är oärlig .
Tom är bedräglig .
Tom är rasande .
Tom är ursinnig .
Tom är gift .
Tom saknas .
Tom är min hjälte .
Tom arbetar .
Tre glassar , tack .
Hon är inte gift .
Han läser allt .
Detta innebar att de var för svaga för att orsaka mer problem .
Han förklarade för min son varför det regnar .
Han var så modig att han inte var rädd för någonting .
Jag hade ingenting att göra med gruppen .
Den här klockan verkar inte fungera som den ska .
Jag läser .
Hans svar är i princip ett nej .
De kommer att komma överens på den punkten .
Han grävde tålmodigt efter fakta .
Länge leve Sovjetunionen !
Hon är upptagen .
Många vet inte om att antibiotika är verkningslösa mot virussjukdomar .
Hon föll ner för stegen .
Välgörenhetsorganisationen har fått sitt namn efter en man som donerade cirka 2 miljarder yen .
Jag har ingen aning om vad jag ska förvänta mig .
Hur går det , sötnos ?
Vilken säng som helst är bättre än ingen säng alls .
Jag glömde att ringa Herr Ford .
Jag skulle vilja ha ett svar .
Det känns som att jag är på bättringsvägen .
Hon ville hjälpa dem .
Lägg köttet i kylen , annars kommer det ruttna .
Han drack direkt från flaskan .
Det är 48 sjömän på skeppet .
Tom har haft problem med sitt vänstra öga sen olyckan .
Jag älskar doften av papper när man slår upp en gammal bok .
Hon är inte ung längre .
Hon är åtminstone 30 år gammal .
Det han sade var inte sant .
Kan du inte ge me lite pengar ?
Har du några syskon ?
Den här typen av smycken har inte mycket värde .
Du luktar så gott .
Jag beordrade ungarna att vara tysta , men de fortstatte att väsnas .
Han pluggar alltid .
Han studerar alltid .
Varför slutar du inte röka ?
Kan någon öppna den här dörren , tack ?
Tom undrade vad Mary ' s efternamn kunde vara .
Glöm inte att signera med ditt namn .
Glöm inte att skriva under med ditt namn .
Det som är svårt att stå ut med är hans överdrivna artighet .
Dykarna hittade ett skeppsvrak på havsbottnen .
Kom igen !
Vi kommer bli sena .
Inga av de här äggen är färska .
Han undvek betet .
Tom låter inte Mary gå och shoppa ensam .
Du borde verkligen sluta röka .
Hennes skämt gick inte hem .
Det här företaget är listat på Parisbörsen .
Mår han bra ?
Han vet hur man flyger en helikopter .
Min son är längre än jag .
I sina böcker rasade han ofta mot regeringen och dess politik .
Jag uppskattar verkligen dina råd .
Får jag lov ?
Han arbetar inte här längre .
Hur står det till ?
Jag har inte sett dig på evigheter !
Han är social av sig .
Festen hölls i professorns ära .
Det regnar idag .
Var är mitt paraply ?
Låt mig betala min del .
Med andra ord : han är lat .
Svaret är helt fel .
Nixon var på väg att bli president .
Tom är förlovad med Ruth .
Reglerna kräver att vi alla är närvarande .
Han kan tala med andar .
Jag kan inte bestämma var vi ska äta lunch ...
Smakar mjölken från den här renen verkligen gott ?
Han tog med henne till vårt ställe .
Var är jag ?
Den här burken är tom.
Hon avskyr honom .
I slutändan är det ändå talangen som räknas i musikens värld .
Jag svettades under armarna .
Tom är inte död .
Tom ser sjuk ut .
Tom ser illamående ut .
Tom saknar dig .
Tom behöver hjälp .
Tom tuppade av .
Tom svimmade .
Tom kolade av .
Tom dog .
Tom verkar trevlig .
Tom kommer inte att stanna .
Vi kan göra det där .
Vi kan inte göra det .
Vi tummade på det .
Vi tog varandra i handen på det .
Vi kommer att vara där .
Vad är de där ?
Vad bryr jag mig om det ?
Hur är den ?
Hurdan är den ?
Hur ser den ut ?
Hur är det ?
Hur känns det ?
Var är de ?
Var är min bil ?
Var är mitt te ?
Vem skulle bry sig ?
Vem håller utkik ?
Vem är på vakt ?
Vem går på vakt ?
Vem är den här killen ?
Vems är de ?
Du kommer att klara dig .
Kan jag få en hund ?
Kan Tom hjälpa oss ?
Missade jag mycket ?
Sa Tom det ?
Sa Tom varför ?
Såg Tom dig ?
Frågade du Tom ?
Varför ge dem någonting ?
Varför frågar du det ?
Varför skulle du fråga det ?
Du kan inte gå ut dit .
Du får inte gå ut dit .
Du kan inte få oss att sluta .
Du kan inte lita på någon .
Du borde inte vara arg .
Du är smartare än jag .
Tyckte du om matchen ?
Hade du roligt på matchen ?
Tyckte du om föreställningen ?
Hade du roligt på föreställningen ?
Tyckte du om rundturen ?
Hade du kul på turnén ?
Tyckte du om rundvandringen ?
Jag luktar med näsan .
Vilka är fördelarna ?
Gjorde du det här ?
Var det du som gjorde det här ?
Hörde du det ?
Såg du Tom ?
Träffade du Tom ?
Använder du droger ?
Tvivlar du på mig ?
Jag är en galning .
Känner du Tom ?
Känner du till Tom ?
Gillar du Tom ?
Tycker du om Tom ?
Älskar du Tom ?
Älskar ni Tom ?
Saknar du Tom ?
Saknar ni Tom ?
Tiden flyger .
Tiden rusar .
Återgå till arbetet .
Hur mår du nu ?
Hur går det ?
Hur är det med Tom ?
Hur går det för Tom ?
Jag kan inte vara säker .
Jag kan inte delta .
Jag kan inte tävla .
Jag kan inte ställa upp .
Jag kan inte göra detta .
Jag kan inte göra det här .
Jag kan inte låtsas .
Jag kan inte bluffa det .
Jag kan inte fejka det .
Jag kan inte hitta den .
Jag kan inte hitta det .
Jag hinner inte .
Jag känner mig illamående .
Jag hatar min röst .
Jag hör skratt .
Jag hörde ett ljud .
Jag hörde ett oljud .
Jag hittade den precis .
Jag hittade det just .
Jag hittade den just .
Jag hittade det precis .
Jag kan allt det här .
Jag vet allt det här .
Jag kan allt detta .
Jag vet allt detta .
Jag gillar din hund .
Jag tycker om din hund .
Jag gillar din hatt .
Jag tycker om din hatt .
Jag älskar det här jobbet .
Jag älskar detta jobb .
Jag älskar detta arbete .
Jag älskar det här arbetet .
Jag älskar er båda .
Jag gjorde den där .
Jag saknar dig , Tom .
Jag behöver en advokat .
Jag behöver dig här .
Jag såg dig aldrig .
Jag såg aldrig dig .
Jag såg aldrig er .
Jag såg er aldrig .
Jag såg Tom i dag .
Jag träffade Tom i dag .
Jag skickade iväg Tom .
Jag skickade hem Tom .
Jag pratade med Tom .
Jag talade med Tom .
Man ska älska sin mamma .
Man ska älska sin mor .
Han tror på det övernaturliga .
Hon väckte honom .
Hon är min typ .
Sitt rakt .
Våren är här .
Våran har kommit .
Den bilen är hans .
Det där är ett bord .
Det där är hans bil .
De är skådespelare .
Vi älskar picknickar .
Vad sa han ?
När kan vi äta ?
Vem är den killen ?
Är du Japansk ?
Är inte du Tom ?
Bob är min kompis .
Kom och hjälp oss .
Var inte arg .
Ställ dig inte upp .
Solen skiner på himlen .
Jag vill ha en advokat .
Jag vill drömma .
Jag önskar dig lycka .
Jag önskar dig allt väl .
Jag önskar dig lycka till .
Jag går och frågar Tom .
Jag ska gå och fråga Tom .
Jag kommer att gå och fråga Tom .
Jag betalar det dubbla .
Jag håller på att bli galen .
Jag blir galen .
Det skulle kunna vara kul .
Det skulle kunna vara roligt .
Det var värt det .
Det är inget problem .
Det är inga problem .
Mary är där inne .
Ni har förändrats .
Jag tror att det är osannolikt att Tom kommer till festen själv .
Tom är ärlig .
Tom är tyst .
Tom har tur .
Tom har anlänt .
Tom är road .
Tom är snabb i vändningarna .
Vi kommer att överleva .
Håll i repet .
Kom när du seger onda drakar , erövrar alla slott och alla prinsessor .
Tom har redan druckit tre koppar kaffe .
Hon äter middag nu .
Tom är säker .
Tom är fortfarande uppe .
Tom är fortfarande vaken .
Det är Tom som bestämmer .
Tom är chef .
Tom är på övervåningen .
Tom är inte glad .
Tom lämnade ett meddelande .
Tom ljög för dig .
Tom ser arg ut .
Tom saknar Mary .
Tom verkade borta .
Tom verkade vilse .
Tom verkade trevlig .
Jag läser ett brev .
Tom bleknade .
Tom blev blek .
Tom var min hjälte .
Tom flämtade .
Tom flåsade .
Tom stönade .
Tom hade helt rätt .
Vänta en sekund .
Vi måste flytta .
Vi måste förflytta oss .
Vad gjorde Tom ?
Vad dödade Tom ?
Vad var det som Tom dödade ?
Vad skrämde dig ?
Jag läste ett brev .
Varför alltid jag ?
Ursäkta mig , talar du engelska ?
Jag älskar Mary så mycket .
Jag vet att ni är upprörda .
Jag vet att du är upprörd .
De är alla oskyldiga barn .
Jag vet att du har rätt .
Jag vet att du mår dåligt .
Jag vet vad som är fel .
Jag vet vad som är rätt .
Jag vet att det är svårt .
Jag vet att detta är svårt .
Jag vet att det här är svårt .
Jag visste att du skulle bli arg .
Jag vill bara prata .
Jag vill bara vila .
Jag hoppas att du har rätt .
Jag hoppas att Tom säger ja .
Jag hörde meddelandet .
Jag har klarsynta drömmar .
Jag har lucida drömmar .
Jag har en annan idé .
Jag hatar att vara dum .
Jag gav Tom ett val .
Jag sov inte bra .
Jag var inte tvungen att åka .
Jag var inte tvungen att gå .
Jag behövde inte åka .
Jag behövde inte gå .
Det fanns ingen där förutom jag .
Det var ingen där förutom jag .
Jag tycker om frukt .
Jag gillar frukt .
Vad fanns inuti ?
Vad heter han ?
Vad finns där inne ?
Vad finns på insidan ?
Vad handlar det om ?
Vad är min belöning ?
Vad är det som är så kul ?
Vad är det som är så roligt ?
Vad är den här till ?
Vad används den här till ?
Vad har du ?
Var är väskan ?
Du babblar .
Du pladdrar .
Du kör så mycket med folk .
Du domderar så mycket .
Du är så kinkig .
Du är så kräsen .
Du kommer med undanflykter .
Är jag i trubbel ?
Är de där till mig ?
Är de där för mig ?
Är de där åt mig ?
Är vi färdiga här ?
Ska vi åka långt ?
Ska vi gå långt ?
Är du en idiot ?
Rodnar du ?
Kan du ta reda på det ?
Kan du se det där ?
Skrev jag det där ?
Sa de hur ?
Sa de varför ?
Blev Tom skadad ?
Skadades Tom ?
Hittade du Tom ?
Hade du roligt ?
Hade du kul ?
Dödade du Tom ?
Kände du Tom ?
Berättade du för Tom ?
Varnade du Tom ?
Klandrar du Tom ?
Förebrår du Tom ?
Lägger du skulden på Tom ?
Litar du på Tom ?
Vill du ha barn ?
Var inte så lat .
Drick inte det där .
Prata inte med mig .
Tala inte med mig .
Berätta inte för någon .
Ha ett bra liv .
Det är bara en tidsfråga .
Tom säger att han aldrig har försökt äta hundmat .
De är alla kannibaler här , utom mig , jag bara blir uppäten .
Båda gick till fönstret för att titta ut .
Min mormor bodde hos oss .
Mannen är naken .
Jag använder Twitter .
Vi är alla överens med er .
Vi är alla överens med dig .
Tom hjälper till .
Du kan ta det .
Du kan ta den .
Jag vek ett hundöra på sidan .
Han är en långväga gäst .
Ibland är det försent att be om ursäkt .
Ha ett trevligt liv .
Allt fungerade problemfritt .
Få Tom att ringa mig .
Han blir rädd lätt .
Han blir lätt rädd .
Han vill ha en iPad .
Hur såg Tom ut ?
Hur visste du ?
Hur ser det ut ?
Hur fungerar det ?
Hur mycket kostar det där ?
Hur mycket är det där ?
Jag kan inte röra det ur fläcken .
Jag kan inte flytta på det .
Jag skulle kunna kyssa dig .
Jag kunde inte stå .
Jag känner inte Tom .
Jag kör en hybrid .
Jag kör en hybridbil .
Jag känner mig så vacker .
Jag blev betalad i dag .
Jag hatar överraskningar .
Jag måste ändra på mig .
Jag hörde det på tv .
Jag hoppas att Tom är okej .
Jag fick precis sparken .
Jag öppnade den precis .
Jag gillar ditt hår .
Jag älskar den sången .
Jag älskar den här delen .
Jag älskar denna del .
Jag älskar den här staden .
Jag älskar denna stad .
Jag älskar dina ögon .
Har du känt honom länge ?
Har du känt henne länge ?
Jag ska resa till Frankrike nästa år .
Det är fullständigt omöjligt .
Desto mer jag tänker på det , desto mindre tycker jag om det .
Han tog expresståget till Tokyo .
Han tog snälltåget till Tokyo .
Jag lär mig språket själv .
Han är inte sjuk .
Han ser trött ut .
Prata inte .
Tala inte .
Le inte .
Vi blir inte yngre .
Vi blir inte yngre än så här .
Tom kom för att hjälpa .
Tom kan höra dig .
Tom kan höra er .
Tom kan inte vägra .
Tom kan inte neka .
Tom kan inte säga nej .
Tom vet inte .
Tom har åkt fast för rattfylleri två gånger .
Tom hjälpte mycket .
Tom är en beatnik .
Tom är en hipster .
Tom är en stamkund .
Tom är en stamgäst .
Tom är fast anställd .
Tom är föräldralös .
Tom är ett föräldralöst barn .
Tom är kompetent .
Tom är skicklig .
Tom är desperat .
Tom ligger i koma .
Tom är eländig .
Tom är olycklig .
Tom är förtvivlad .
Tom är för ung .
Tom gillar det hett .
Tom gillar det varmt .
Tom gillar den varm .
Tom såg bra ut .
Tom ser skyldig ut .
Tom vill ha en kyss .
Tom vill ha en puss .
Tom blev kidnappad .
Tom blev bortförd .
Tom blev bortrövad .
Jag blev bortförd av utomjordingar .
Jag blev bortförd av rymdvarelser .
Jag blev kidnappad av rymdvarelser .
Jag blev kidnappad av utomjordingar .
Enlevering är en så gott som utdöd företeelse i Sverige .
Nuförtiden är sms-avisering lika vanligt som brevavisering .
Här är bussen .
Vilken är din favoritsuperhjälte ?
Vem är din favoritsuperhjälte ?
Jag litar på dig .
Tom är smart .
Det ligger tre grytunderlägg på bordet .
Är det några frågor ?
Tom har åkt .
Tom är borta .
Tom är fri .
Tom är tjock .
Tom är full .
Tom blev arresterad .
Tom lyssnar inte .
Blev Tom mördad ?
Det kan vi inte göra .
Vi måste skynda oss .
Blev du beskjuten ?
Vad sa Tom ?
Vad missade vi ?
Vad träffade du ?
Vad såg du ?
Vad vet du ?
Vad är allt det här ?
Vad är allt detta ?
Vad är det här för ?
Vad är det här till ?
Vad är detta för ?
Vad är detta till ?
Vadan denna panik ?
Vad har Tom hittat ?
Vad är din plan ?
Vad är er plan ?
Vad har du gjort ?
Vad har ni gjort ?
När börjar vi ?
När startar vi ?
Var är vi nu ?
Vart gick Tom ?
Var är alla ?
Var är allihopa ?
Var är allesammans ?
Var är min telefon ?
Varför är du hemma ?
Varför är ni hemma ?
Vi har problem .
Vi är i trubbel .
Vi är illa ute .
Vi är i knipa .
Vi har råkat illa ut .
Ska du ut ?
Kan jag få prata med dig ?
Kan Tom få en hund ?
Sa de när ?
Kom Tom tillbaka ?
Hans dumma svar överraskade allihopa .
Hans dumma svar överraskade alla .
Herr White är en förnuftets man .
Herr White är en förnuftig man .
Hon är orolig över din säkerhet .
Hon är orolig över er säkerhet .
Vi är benägna att slösa tid .
Jag läser spanska .
Jag studerar spanska .
Jag trodde att det skulle vara värt det .
Jag tänkte att det skulle vara värt det .
Var är satelliterna ?
Tom gillar inte Marys attityd .
Tom tycker inte om Marys attityd .
Kysste du Mary ?
Pussade du Mary ?
Vill du ha ett jobb ?
Vill du ha ett arbete ?
Vet Tom än ?
Rör inte dem .
Tycker du inte om mig ?
Har Tom blivit skadad ?
Har Tom skadats ?
Har du sett Tom ?
Hennes dröm är över .
Hennes hud var varm .
Hur illa kan det vara ?
Hur dåligt kan det vara ?
Hur dålig kan den vara ?
Flodens övre lopp är mycket vackert .
Vad är det för fel på honom ?
Hon dog av törst under torkan .
Hur gissade du ?
Hur kunde du gissa ?
Hur klarar du det ?
Hur lyckas du ?
Jag uppskattar det .
Jag kan inte förneka det .
Jag kan inte behålla det här .
Jag kan inte behålla den här .
Jag kan inte lämna dig .
Jag kunde inte säga nej .
Jag gjorde dig en tjänst .
Jag dödade inte Tom .
Jag känner mig inte sjuk .
Jag vill inte ha det här .
Jag vill inte ha den här .
Jag vill inte ha denna .
Jag vill inte ha detta .
Jag måste få träffa Tom .
Jag måste träffa Tom .
Jag har arbete att göra .
Jag vet bara inte .
Jag vet vem som gjorde det .
Jag gillar att vara upptagen .
Jag gillar den där tröjan .
Jag gillar den där skjortan .
Jag gillar din scarf .
Jag gillar din halsduk .
Jag gillar din sjal .
Jag gillar din sjalett .
Jag tycker om din scarf .
Jag tycker om din halsduk .
Jag tycker om din sjal .
Jag tycker om din sjalett .
Ljuger du för mig ?
Vi har varit uppe hela natten .
Jag tappade ett örhänge .
Jag älskar den där klänningen .
Jag älskar den filmen .
Jag älskar den scarfen .
Jag älskar den halsduken .
Jag älskar den sjalen .
Jag älskar den sjaletten .
Jag älskar den berättelsen .
Jag älskar den historian .
Jag älskar den sagan .
Jag behöver en huvudvärkstablett .
Jag behöver lite sömn .
Jag behöver lite vatten .
Jag behöver få träffa Tom .
Jag behöver träffa Tom .
Nej , inte riktigt .
Hon sprang så fort som hon förmådde .
Amerika är ett land av invandrare .
Gott Nytt År !
Tom backade inte ut .
Tom sprang efter Mary .
Jag räddade ditt liv .
Jag träffade Tom i kväll .
Jag såg Tom i kväll .
Jag förstår vad problemet är .
Jag vill vara här .
Jag vill åka tillbaka .
Jag vill gå tillbaka .
Jag vill träffa Tom .
Jag var på området .
Jag hämtar lite is .
Jag hämtar boken .
Jag ska hämta boken .
Jag undersöka det .
Jag forska i det .
Jag ska jobba på det .
Jag är lite upptagen .
Jag är en tålmodig man .
Jag är alldeles ensam nu .
Jag är helt ensam nu .
Jag är hemskt trött .
Jag kommer till dig .
Jag ska skaffa katt .
Jag är glad att vi är överens .
Jag chansar bara .
Jag är precis som du .
Jag är sen till jobbet .
Jag är sen till arbetet .
Jag ger inte upp .
Det är svårt att säga .
Låt oss göra affärer .
Har den ett badrum ?
Var tålmodig .
Ha tålamod .
Var tålmodiga .
Han blev ditsatt för mord .
Han blev falskeligen anklagad för mord .
Han blev snärjd för mord .
Vart gick han ?
Vi sätter julgranen här .
Vi ställer julgranen här .
Lägenhet är försedd med både förråd och balkong .
Divanen är en populär soffmodell .
I Grekland förvärras skuldkrisen .
Seoul är huvudstaden i Sydkorea .
Han dog innan jag kommit fram .
Han dog innan jag kom fram .
Överlappning kan inträffa .
Underteckna på den här raden .
Signera på raden här .
Sluta trakassera mig .
Sluta besvära mig .
Berätta för mig om Tom .
Det var poängen .
De är dyra .
Detta är inkorrekt .
Det här är inkorrekt .
Detta är oriktigt .
Det här är oriktigt .
Detta är felaktigt .
Det här är felaktigt .
Så kan Tom inte göra .
Tom kan inte göra så .
Tom kan inte göra det .
Tom får inte göra det .
Tom kan inte skada mig .
Tom får inte skada mig .
Tom kan inte se dig .
Tom får inte se dig .
Tom kan inte träffa dig .
Tom får inte träffa dig .
Tom såg det inte .
Tom såg inte det .
Tom hade inget val .
Tom är skadad .
Tom har blivit skadad .
Tom skadade knät .
Tom är en korgosse .
Tom är sångare i gosskör .
Tom är en flykting .
Tom är en rymling .
Tom är en landsflykting .
Tom är på baren .
Tom är bakom dig .
Tom är illa ute .
Tom är i knipa .
Tom har problem .
Tom är min make .
Tom är min man .
Helsingfors är Finlands huvudstad .
Tom kommer inte .
Tom är på väg .
Tom är otrogen .
Tom är trolös .
Tom är klarvaken .
Tom sitter inte i fängelse .
Tom är inte i häkte .
Tom sitter inte i häkte .
Tom gillar det kallt .
Tom ser irriterad ut .
Tom ser besvärad ut .
Tom ser förkrossad ut .
Tom behöver en tjänst .
Tom lurade mig .
Tom såg videon .
Om du inte studerar mer så kommer du helt säkert att misslyckas .
Hon kom in helt tårögd .
Endast då förstod jag vad han menade .
Jag kan inte se något med mitt högra öga .
Jag oroar mig inte så mycket om mitt CV .
Detta är hyddan som han levde i .
Jag såg en gammal vän .
Hunden är på stolen .
Mary har många vänner .
Jag har köpt en bil .
Jag har inte råd att betala så mycket .
Släpp henne .
Bess är endast ett barn .
Kan du inte skriva " Pfirsichbäumchen " ?
Det är så simpelt .
Kan du hålla det en hemlighet ?
Var snäll och påminn mig om jag glömmer bort .
Ingen visste att du var i Tyskland .
En katt är inte en person .
Den här ordboken kan komma till användning .
Hon gillade poesi och musik .
Har du namngett din nyfödda bäbis ?
Jag är inte din slav .
De vill inte att du ska veta .
Tom tackade Mary för hennes råd .
Tom vet Marys hunds namn .
Hans uppfinning är överlägsen konventionell utrustning .
Hur många självmord tror du att det sker varje år i Japan ?
Du hade läst .
Sluta upp med det omedelbart .
Han är bara en amatör .
Du borde inte titta ner på honom .
Å ena sidan är han snäll men å andra sidan är han lat .
Vi föddes på samma dag .
Fem gånger sju är trettiofem .
Det verkar som att han känner till det .
När kan vi mötas igen ?
" Det är första gången jag river min ägare " , sa katten .
Tom fick inte något gjort idag .
Ju mer du lär känna henne , desto mer kommer du att gilla henne .
Jag tyckte jag sa åt dig att inte stå i vägen för mig .
Var finns närmaste hotell ?
Tom skrattade sällan åt Marys skämt .
Schweiz är beläget mellan Frankrike , Italien , Österrike och Tyskland .
Jag trodde att du hade en överenskommelse med Tom .
Hon sa att hon hade en förkylning .
Vi insåg inte att vi var så högljudda .
Jag vill ha en massage .
Jag behöver slappna av .
Vi kan inte ge upp utan en kamp .
Mor , far .
Titta på ert lilla monster .
Min dröm är att leva fredfullt i byn .
Han slåss mot väderkvarnar .
Tom frågade Mary om hon kunde hjälpa honom .
Kommer du ihåg oss ?
Hon väntar .
Du har många vänner .
Hon valde en hatt som matchade hennes klänning .
Det här klassrummet är städat .
Det var fönstret som Jack tog sönder igår .
Vi är bekanta med den här sången .
Är din lägenhet väl underhållen ?
Du älskar kaffe .
Tom tycker inte om huset han bor i .
Vi sover vanligtvis i det här rummet .
De som styr mest gör minst ljud ifrån sig .
Detta är en kamera tillverkad i Japan .
Var är tvättrummet ?
På grund av den dåliga skörden har vetepriset gått upp de senaste sex månaderna .
Jag var oförmögen att titta henne i ansiktet .
Kaffet var så varmt så jag inte kunde dricka det .
Kan du visa mig en billigare kamera än denna ?
Kan jag få ett glas vatten , tack .
Tom säger att han är villig att göra det gratis .
Jag kan inte gå förrän han kommer .
Vår värd erbjöd oss en drink .
Massorna reste sig mot diktatorn .
Allt var fortfarande i skogen .
Håll repet .
Kan du vakta ungarna ?
Hittade dom någonting ?
Vann du trofén ?
Vet du vem han var ?
Blir du ledsen av det ?
Vet Tom vem jag är ?
Ser Tom förvirrad ut ?
Smickra inte dig själv .
Lova att du inte blir arg .
Gå inte ut på framsidan .
Få mig inte att skada dig .
Få mig inte att döda dig .
Slösa inte bort Toms tid .
Oroa dig inte .
Det är enkelt .
Tar du dörren ?
Få bort Tom härifrån .
Gå hem .
Vila upp dig .
Han är mörk och snygg .
Hur mycket kostade det ?
Jag uppskattar din tid .
Jag uppskattar ditt jobb .
Jag kan inte komma just nu .
Jag kan inte hantera det här .
Vad tycker du om den här tröjan ?
Det här är den vackraste blomman i trädgården .
Tom brukade hata Mary .
Nu älskar han henne .
Du borde ha kommit med oss .
Den första gruppen studerar på morgonen , den andra på kvällen .
Ut härifrån !
Allihopa !
Till och med en bra dator kan inte klå dig på schack .
Vi visste inte vad vi skulle göra .
Vi kysstes bara .
Tom tycker att det är tillräckligt bra .
Jag sa inte att det inte var okej att äta .
Många människor litar inte på regeringen .
Katten sover på soffan .
Hon köpte en bok i affären .
Vem tycker inte så ?
Jag hoppas att du njuter av din vistelse här .
Jag kommer tillbaka om 2 veckor .
Jag har så mycket arbete så jag stannar en timme till .
Han skyndade sig tillbaka från England .
Jag känner mig väldigt kall .
Peter är inte alls lik hans pappa .
Låt oss hoppas på bra resultat .
Han sparkade honom medan han låg ner .
Tom gjorde ett halv-färdigt jobb .
Jag föddes här .
Träning är för kroppen , vad läsning är för sinnet .
Huset brann ner till grunden .
Tom håller på att somna .
Han är duktig med kort .
Bonde plöjde hans fält hela dagen .
Du behöver inte vänta till slutet .
Hon kände sig illa till mods vid tanken på hennes framtid .
Det var en tyst natt i vintertid .
Tårta ?
Jag blev plötsligt hungrig igen .
Förlusten av hennes far var väldigt smärtsamt för henne .
Alla studenterna i klassen gillar herr Smith .
Jag vinkade av honom vid flygplatsen .
Vilken nagellack är din favorit ?
Skeppet sjunker .
Tycker du om teatern ?
Du borde lita på mig .
Mary har redan gått .
En liten vinst är bättre än en stor förlust .
Hon dog 1960 .
Jag brukade simma i havet när jag var ett barn .
Jag hade en intressant konversation med min granne .
Tom förlät Mary på hennes dödsbädd .
Det råder ingen tvekan om att hon älskar honom , men hon vill inte gifta sig med honom .
Livet är ett uppvaknande efter ett annat .
Gå och byt om .
Mohand är min halvbror .
Det fanns lite dagg imorse .
Detta är min lärare .
Han heter herr Haddad .
Hans hobby är att samla på gamla frimärken .
Hur många århundraden finns det på ett millennium ?
Han var rädd att du skulle skjuta honom .
Var skulle du vilja åka nästa söndag ?
Har du en kofot i verktygslådan ?
Livet är inte lätt .
Hon övergav sina barn .
Nej , inte för mycket .
Ditt svar på frågan visade sig vara fel .
Jag förstod inte hans skämt .
Har du borstat tänderna ?
Mary ser ovänlig ut , men egentligen har hon ett gott hjärta .
Jag kände ett tryck på min axel och vände mig om .
Jag är egentligen en universitetslärare .
Det är tystnad som är dyrbart nu .
Jag är så stolt över dig .
Att lära sig koreanska är svårt .
Kan du släppa av mig vid biblioteket ?
Jag har beslutat mig för att svara på alla frågor offentligt .
Katten flydde med en bit fisk från köket .
Katten klängde vid hennes klänning .
Kvinnor känner att män ofta är väldigt komplicerade .
Min mamma lagar mat åt mig .
Tom ville hämnas .
Jag träffade honom en gång .
Franskan utvecklades från latin .
Väggarna i det gamla huset var inte raka .
Han må vara ung , men han är verkligen en tillförlitlig person .
Det är inte nödvändigt för oss att närvara vid mötet .
Den mänskliga handen har fem fingrar med naglar .
Den nya telefonboken är här !
Spara lite glass åt mig .
Vi är femton , allt som allt .
Jag har inte sett henne sen förra månaden .
Jag skulle vilja byta rum .
Min bror är lika lång som jag .
Bilal är utbildad .
Jag tror att jag äntligen ska pensionera mig .
Hon var tvungen att ge upp planen .
Hon har tagit på sig alltför mycket arbete .
Han bröt nacken i olyckan .
Han kände sig obekväm i hans fars närvaro .
Kate låg ner med öppna ögon .
Roy behövde inte skynda sig till flygplatsen för att möta hans föräldrar .
Han löste korsordet med lätthet .
Jag har fortfarande inte funnit det jag söker efter .
Jag har fortfarande inte hittat det jag letar efter .
Hans historia är sann .
Ett högt träd kastar sin långa skugga på vattnet .
Var god , kryssa i den lämpliga rutan .
Han ska övertala sin far att köpa en ny bil .
Hon går ofta och shoppar på helger .
Det dröjer inte länge innan hon är tillbaka .
Du kan komma och se mig närhelst det passar dig .
Ge mig en till kopp kaffe .
Är det säkert att simma i den här floden ?
Jag ville träffa dig .
Jag kunde svära på att någonting rörde sig .
Om jag var rik så skulle jag åka utomlands .
Tom visste att jag var på väg .
Det var ett väldigt spännande spel .
Hon kommer att betala för allting .
Jag önskar att jag hade en bil .
Stanna gärna kvar efter konserten .
Vi kommer signera autografer .
Jag är älskad av mina föräldrar .
Är du för eller emot planen ?
Jag gick också .
Jag menade inte något av det .
Jag uppskattar verkligen din hjälp .
Av någon anledning så känner jag mig mer levande på natten .
Jag vill bara ha roligt .
Vad är det med dig ?
Tom vill ha hjälp .
Tom vill leka .
Tom vill spela .
Tom var deprimerad .
Tom kommer att vara här .
Titta på hur jag gör det .
Titta hur jag gör det .
Vad gör vi ?
Kolla hur jag gör det .
Vad visste Tom ?
Vad ville Tom ?
Vad ville Tom ha ?
Vad gör jag härnäst ?
Vad gör jag sen ?
Vad är jag skyldig dig ?
Vad är jag skyldig er ?
Glad mors dag !
Vad gör vi nu ?
Vad är det som luktar ?
Vad är det där för lukt ?
Stör jag dig ?
Middagen var toppen .
Tycker du om robotar ?
Behöver du en hand ?
Var inte arg på mig .
Bli inte paranoid .
Släpp mig inte .
Släpp inte taget om mig .
Ställ inte till en scen .
Tacka mig inte än .
Se till att Tom ringer mig .
Ge Tom allting .
Gå och hämta lite handdukar .
Gå och vänta i bilen .
Har du sett det här ?
Han föste iväg henne .
Han är en drama queen .
Hon är en drama queen .
Hur kan vi göra det ?
Hur kom Tom in ?
Hur tog sig Tom in ?
Hur tog Tom sig in ?
Hur känns det där ?
Jag tror att Tom ljög för oss .
Någon måste vara här för barnen .
Hon förlorade sina pengar , sin familj och sina vänner .
Det gläder mig att höra om den nyfödde .
Det glädjer mig att höra om den nyfödde .
Han gladdes av sällskapet .
Skulle du kunna förklara vägen till Madame Tussaud ?
Skulle ni kunna förklara vägen till Madame Tussaud ?
Bara kärlek kan krossa ditt hjärta .
Bara kärlek kan krossa hjärtat .
Bara kärlek kan krossa ens hjärta .
Endast kärlek kan krossa ditt hjärta .
Endast kärlek kan krossa hjärtat .
Endast kärlek kan krossa ens hjärta .
Nu är hon precis fyra .
Staden förstördes under kriget .
Varför frågar du inte din lärare om råd ?
Han är alltid full av livskraft .
Han är alltid full av energi .
Han är alltid en man vid full vigör .
Min engelska är allt men inte bra .
Min engelska är allt utom bra .
Min engelska är inte alls bra .
Tom är inte en bra kock .
Jag har försökt att lösa det här problemet i timmar .
Hur ser det här ut ?
Hur svårt kan det vara ?
Hur skulle du veta ?
Hur kom du hit ?
Hur tog du dig hit ?
Hur mår du ?
Hur känner du dig ?
Hur mår din patient ?
Jag kan höra vinden .
Jag kan inte tillåta det .
Jag kan inte bryta mig loss .
Jag kan inte bryta mig fri .
Jag kan inte bekräfta det .
Jag lånade honom lite pengar , men han har inte betalat tillbaka dem än .
Jag lånade honom lite pengar , men har inte återbetalat dem än .
Jag tar det som ett tecken på kärlek .
Jag tål inte golf .
Jag dubbelkollade det .
Jag kollade det två gånger .
Jag kontrollerade det två gånger .
Jag gjorde det frivilligt .
Jag rörde inte Tom .
Jag ville inte ha mjölk .
Jag kände mig skyldig .
Jag hittade din dagbok .
Jag måste åka hem .
Jag måste ta mig hem .
Jag hoppas att vi hittar Tom .
Jag fann din dagbok .
Jag hoppas att vi finner Tom .
Konstiga saker hände på hennes födelsedag .
Konstiga saker skedde på hennes födelsedag .
" Vad tänker du på ? "
" Jag tänker på dig . "
Romanen är mycket rörande .
Vi kommer ifrån olika länder .
Har du sett Shaoxingopera ?
Han är alltid kvick och slagfärdig .
Hon hade ett litet , runt föremål i handen .
Han hade ett litet , runt föremål i handen .
Ät den här .
Ät det här .
Ät denna .
Ät detta .
Jag är less på att vara pensionerad .
Jag är trött på att vara pensionerad .
Hon gav mig inte sitt namn .
Det är ett rökmoln över landskapet .
Det är ett rökmoln över provinsen .
Jag lånade den precis .
Jag lånade den bara .
Jag kan bara inte sova .
Jag kan inte sova bara .
Jag ville bara ha pengar .
Jag kände din far .
Jag kände din fader .
Jag kände din pappa .
Jag vet vad jag vill .
Jag vet vad jag vill ha .
Jag vet att du är upptagen .
Jag vet att ni är upptagna .
Jag gillade den där filmen .
Jag gillade den filmen .
Jag gillade din historia .
Jag tyckte om din historia .
Jag älskar utmaningar .
Jag saknar Tom så mycket .
Jag rörde den aldrig .
Jag läste din rapport .
Jag såg vad Tom gjorde .
Jag såg vad du gjorde .
Jag tror att jag gillar dig .
Jag trodde att du slutade .
Jag trodde att du slutat .
Jag var ironisk .
Jag var artig .
Jag var hövlig .
Han visade mig massor av vackra bilder .
Jag skulle vilja träffa Tom .
Jag är lite tidig .
Jag är fotograf .
Jag är lealös .
Jag är mjuk i lederna som en akrobat .
Det har blivit märkbart kallare .
Tror du att Steve Jobs skulle ha varit lika framgångsrik som han varit om hans efternamn varit " Joobs " istället ?
Om du inte vill att jag ska åka , så gör jag det inte .
Vissa studenter kommer inte att komma tillbaka nästa termin .
Några studenter kommer inte att komma tillbaka nästa termin .
Han vred om min arm .
Han utövade påtryckningar på mig .
Tom hjälper .
Var kan jag köpa frimärken ?
Skulle du kunna sänka radion ?
Tom är egensinnig .
Vi flög från London till New York .
Hon liknar inte sin mor alls .
Hon liknar inte inte sin mamma alls .
Smickrare liknar vänner , på samma sätt som vargar liknar hundar .
Smickrare liknar vänner , liksom vargar liknar hundar .
Vi liknar verkligen inte varandra .
En fladdermus som flyger på himlen liknar en fjäril .
Om du anstränger dig kan du förbättra din engelska .
Enligt tidningen begick han självmord .
Jag skulle vilja gå och sova nu .
Den är två gånger så stor som denna .
Den är dubbelt så stor som denna .
Kommittén sammanträder två gånger om månaden .
Kommittén sammanträder två gånger i månaden .
Kommittén sammanträder två gånger per månad .
Ja !
Jag vann två gånger i rad .
Vi väntade .
Han kommer att komma .
Här kommer Tom .
Vad du har växt !
Tjejer kom in , den ena efter den andra .
Flickor kom in , den ena efter den andra .
Vet du vem Rie Miyazawa är ?
Han stannade där hela tiden .
Jag tog Tom till sjukhuset .
Hur länge ska du vara i Japan ?
Jag känner mig hungrig .
Jag håller på att bli bättre .
Jag följer med Tom .
Jag är så generad .
Det slutade bra .
Det var mitt nöje .
Släng iväg den bara .
Kasta den bara .
Ur vägen för mig .
Håll dig ur min väg .
Håll er ur min väg .
Oroa dig inte .
Han förstår inte tyska .
Oroa dig inte .
Han kan inte tyska .
Alice sover i mitt rum .
Låt mig hjälpa dig upp .
Låt mig prata med Tom .
Låt mig tala med Tom .
Mina väskor är packade .
Återvänd till skeppet .
Så vad gjorde du ?
Håll dig borta från Tom .
Stanna här med Tom .
Stanna , annars skjuter jag .
Sluta prata med mig .
Hälsa till Tom .
Hälsa Tom att jag är färdig .
Säg till Tom att jag är färdig .
Det där är ett gammalt skämt .
Detta är skandalöst !
Det här är skandalöst !
Det här är riktigt illa .
Detta är riktigt illa .
Det här är väldigt färskt .
Det här är inte korrekt .
Det här är inte riktigt .
Tom åt upp ditt godis .
Tom spelar på hästar .
Tom är sannerligen en mångsysslare .
Tom har många dåliga vanor .
Tom ger upphov till betydligt många fler meningar än Mary .
Jag gillar inte att bli driven med .
Det här problemet är för svårt att lösa för lågstadieelever .
Jag lagar kyckling .
Det här arbetet är inte på något sätt lätt .
Tom sjukanmälde sig .
Tom hör dig inte .
Tom kan inte höra dig .
Tom kan inte skada dig .
Tom skulle kunna vara en polis .
Tom berättade inte det för mig .
Tom äter som en gris .
Tom satte sig i bilen .
Tom har svimmat .
Tom har tuppat av .
Tom har kolat av .
Tom måste gå hem .
Tom är en bra grabb .
Du måste inte bestämma dig just nu .
Hur mår din mor ?
Hur mår din mamma ?
Jag heter Henry .
Du måste lämna Boston .
Han kommer alltid att älska henne .
Varför behöver du de här pengarna ?
Varför behöver du dessa pengar ?
Vad tycker du om att göra på söndagar ?
Vad gillar du att göra på söndagar ?
Det är någonting med honom som jag inte tycker om .
Jag tycker att du är lite för försiktig .
Jag tror att du är lite för försiktig .
Jag tycker att du är lite för noggrann .
Jag tror att du är lite för noggrann .
Allt måste handskas med väldigt försiktigt .
Du borde vara försiktigare nästa gång .
Du borde vara noggrannare nästa gång .
Ni borde vara försiktigare nästa gång .
Ni borde vara noggrannare nästa gång .
Tom är en smart grabb .
Tom är sociopat .
Tom ska precis gå .
Tom är vid dörren .
Tom kommer tillbaka .
Tom är mållös .
Tom är förbluffad .
Tom är häpen .
Tom är förstummad .
Tom har aldrig fel .
Tom är på lastkajen .
Tom är på lastningsplatsen .
Tom är precis här .
Tom är här .
Tom är fortfarande vid liv .
Tom är omöjlig att hindra .
Tom är omöjlig att stoppa .
Tom är ohejdbar .
Tom dök precis upp .
Tom dök bara upp .
Tom var medveten om riskerna .
Tom tittade på Mary .
Tom såg förbryllad ut .
Tom såg villrådig ut .
Tom såg häpen ut .
Tom såg frågande ut .
Tom ser orolig ut .
Tom ser upphetsad ut .
Tom ser upprörd ut .
Tom ser förvirrad ut .
Tom ser konfys ut .
Tom ser konfunderad ut .
Tom ser omtumlad ut .
Jorden är där vi alla bor .
Jordens latinska namn är Tellus .
Jordens namn på latin är Tellus .
Jag trodde att ni två var lika gamla .
Han glömmer aldrig att skicka en födelsedagspresent till sin mor .
Han glömmer aldrig att skicka en födelsedagspresent till sin mamma .
Flera i partitoppen har fått avgå .
Kärleken är till sin natur blind .
Jag behöver en askkopp .
Han undersökte Amazonas regnskog .
Han utforskade Amazonas regnskog .
Han genomforskade Amazonas regnskog .
Vad är det som du säger ?
Tom ser bekant ut .
Tom ser ut som du .
Tom ser lättad ut .
Tom fick Mary att sluta .
Tom har kanske rätt .
Tom måste hjälpas .
Tom måste få hjälp .
Tom verkar stressad .
Tom skickade mig ett meddelande .
Tom skakade på huvudet .
Tom borde vara här .
Tom var otrolig .
Tom var ofattbar .
Tom var fantastisk .
Tom var väldigt modig .
Tom skrek åt Mary .
Tom skrek på Mary .
Blev någon dödad ?
Vi kan inte dödas .
Vi får inte dödas .
Vi kan inte göra det nu .
Vi får inte göra det nu .
Vi har inga hemligheter .
Vi borde ringa Tom .
Vi klarar oss .
Vi kommer att klara oss .
Vi har pratat färdigt .
Vi kommer att försöka .
Vi är sena .
Stod ni två nära varandra ?
Vad ville de ?
Vad lärde du dig ?
Vad hände sen ?
Vilken station är det här ?
Vilken station är detta ?
Vad skulle ha veta ?
Varför dröjer Tom ?
Vad uppehåller Tom ?
Vad är avbrottet ?
Du äter inte någonting .
Vad är det med Tom ?
När kommer Tom ?
När är begravningen ?
Du kan inte backa ur .
Du får inte backa ur .
Du kan inte hoppa av .
Du får inte hoppa av .
Du får inte smita .
Du kan inte skylla på mig .
Du får inte skylla på mig .
Du får inte ringa Tom .
Du får inte skada Tom .
Du kan inte skada Tom .
Ni får inte skada Tom .
Ni kan inte skada Tom .
Var bodde du ?
Var bodde ni ?
Han dricker inte .
Du kan inte lämna mig .
Du får inte lämna mig .
Ni kan inte lämna mig .
Ni får inte lämna mig .
Du kan inte sluta nu .
Du får inte sluta nu .
Ni får inte sluta nu .
Ni kan inte sluta nu .
Du hjälper inte till .
Ni hjälper inte till .
Du är så paranoid .
Ni är så paranoida .
Tyckte du om det där ?
Njöt du av det där ?
Stör jag er ?
Är du polis ?
Är du polisman ?
Kan vi bara gå hem ?
Kom och träffa allihop .
Berättade någon för Tom ?
Förlät Tom dig ?
Har du gått ned i vikt ?
Har vi något val ?
Behöver vi en plan B ?
Har du en telefon ?
Har ni en telefon ?
Ser du någonting ?
Ser ni någonting ?
Spela inte förvånad .
Avbryt inte Tom .
Han vände bort blicken .
Han festar för mycket .
Hans föräldrar älskar mig .
Den här bilen är inte lika fin som den där .
Hur kan vi rädda Tom ?
Hur hände det där ?
Hur hittade Tom oss ?
Hur hittade ni oss ?
Hur hittade du oss ?
Hur känner du Tom ?
Hur känner ni Tom ?
Hur länge har vi på oss ?
Hur lång tid har vi ?
Hur ska du klara dig ?
Hur ska ni klara er ?
Jag kan inte svara på det .
Jag kan inte ändra på det .
Jag kan inte kontakta Tom .
Jag får inte kontakt med Tom .
Jag kan inte få kontakt med Tom .
Jag kan inte kontrollera Tom .
Jag kan inte göra mer .
Jag kan inte göra det själv .
Jag klarar det inte själv .
Jag kan inte göra det i dag .
Jag klarar det inte i dag .
Jag kan inte göra det nu .
Jag klara det inte nu .
Jag kan inte rita en fågel .
Jag kan inte titta på Tom .
Jag klarar inte av lögnare .
Jag står inte ut med lögnare .
Det kommer antagligen att snöa i morgon .
Det där var riktigt kul .
Gör det igen !
Det där var riktigt roligt .
Gör det igen !
Läs detta först .
Läs det här först .
Jag vill inte träffa någon i dag .
Jag börjar komma ihåg det .
Det här nyttar ingen .
Det där är i hög grad en viljesak .
Jag kanske kommer att prata med Tom .
Jag kanske pratar med Tom .
Jag behöver bilnycklarna .
Jag rörde aldrig Tom .
Jag träffar Tom varje dag .
Jag ser Tom varje dag .
Jag borde inte vara här .
Jag stal den från Tom .
Jag stal det från Tom .
Jag tror att jag är förälskad .
Jag tror att jag är kär .
Jag tycker att du är trevlig .
Jag tycker att du är snäll .
Jag tänkte på Tom .
Jag sa åt dig att gå .
Jag sa åt er att gå .
Jag sa åt dig att ge dig iväg .
Jag sa åt er att ge er iväg .
Jag försökte varna dig .
Jag försökte varna er .
Jag vill be om ursäkt .
Jag vill komma hem .
Jag skulle dö utan dig .
Jag skulle dö utan er .
Jag skulle vilja se Tom .
Jag ringer efter en taxi åt dig .
Jag ringer en taxi åt dig .
Jag betalar på mitt eget sätt .
Jag berättar för Tom senare .
Jag ska berätta för Tom senare .
Tusen tack för din vänlighet .
Tusen tack för er vänlighet .
Tack för ditt svar .
Tack för ert svar .
Vi är tacksamma för er vänlighet .
Vi är tacksamma för din vänlighet .
Ett stort tack för din hjälp .
Ett stort tack för er hjälp .
Tack för er gästfrihet .
Tack för din gästfrihet .
Tack för ditt hårda arbete .
Tack för ert hårda arbete .
Var ska vi träffas ?
Var ska vi ses ?
Härifrån till banken är det gott och väl tre kilometer .
Jag är socialarbetare .
Jag är oskyldig .
Jag är en oskyldig man .
Jag ska gå nu .
Jag kommer att gå nu .
Jag går nu .
Det hände så snabbt .
Det var bara en liten kärleksaffär .
Det var fortfarande riktigt varmt , trots att solen hade sjunkit ganska lågt .
Följ efter bilen .
Jag har varit bekant med henne i över 20 år .
Jag har känt henne i över 20 år .
Jag ser .
Klä på er .
Hitta Tom .
Stå inte .
Skrik inte .
Han nämnde det .
Vilken tand gör ont ?
Tom är stark .
Tom är sträng .
Tom är blyg .
Tom är ledsen .
Tom har rätt .
Det är kvavt här inne .
Det är kvalmigt här inne .
John fick Mary att hoppa till .
John fick Mary att hoppa .
Berätta bara inte för Tom .
Följ bara mitt exempel .
Mary är ganska orolig .
Mary är ganska stökig .
Någon satte dit honom .
Stanna där du är !
Stanna där ni är !
Sluta kalla mig för Tom .
Sluta anmärka på Tom .
Sluta hacka på Tom .
Säg till Tom att jag älskar honom .
Berätta för Tom att jag älskar honom .
Det står en man med en pistol i handen i dörren .
Det står en man med en pistol i handen vid dörren .
Rökning är skadligt .
Vi gör mjölk till ost och smör .
Vi gör ost och smör av mjölk .
Tom har gått .
Tom är glad .
Tom är snabb .
Tom har dött .
Det såg billigt ut .
Det är lunchdags .
Är det vitt ?
Jag bor här .
Jag gillar te .
Vi förlorade .
Det var en bra dag .
Hon sprang så fort hon kunde .
Nöden är uppfinningarnas moder .
Turkisk lira är den officiella valutan i Turkiet .
Jag är galen .
Jag är ledsen , men jag har ingen växel .
Han var beredd att ge tillbaka till henne alla hennes pengar .
Ring till polisstationen och berätta för dem vad du berättade för mig .
Idén var så avancerad att jag inte förstod den .
Kyckling , tack .
Tom la på telefonen .
Tom lade på telefonen .
Tom drog sig inte ur .
Tom tänkte inte tillbaka .
Tom skulle kunna vara var som helst .
Tom åt en snabblunch .
Tom åt en snabb lunch .
Vi kommer att vinna .
Lova mig att du inte berättar för henne .
Tom högg tag i sin väska .
Tom grep tag i sin väska .
Tom ryckte till sig sin väska .
Tom höll Mary tätt .
Tom hjälpte oss mycket .
Tom la på i örat på Mary .
Tom är tillbaka i stan .
Tom är knappt vid liv .
Tom är besviken .
Tom skalade potatis .
Tom ignorerar dig .
Tom är uppe på vinden .
Tom sover fortfarande .
Tom gråter fortfarande .
Tom är deras ledare .
Tom är för långt borta .
Tom andas inte .
Det är inte Tom som bestämmer .
Vi ska vinna .
Tom är farlig .
Strävan efter sanning är beundransvärd .
Ha det så kul !
Hur så ?
Jag vill lära mig lettiska .
Å , det är en världslig sak !
Varsågod att ta plats !
Var god och ta plats !
Han vill inte att du berättar för honom om ditt sexliv .
Han vill inte att du berättar för honom om ert sexliv .
Han vill inte att ni berättar för honom om ert sexliv .
Snälla prata inte så snabbt .
Vänligen , prata inte så snabbt .
Jag borde sluta skjuta upp saker och ting .
Kyrkan är mitt i byn .
Han kommer att gå .
Tom går till skolan till fots .
Livet i fängelse är värre än ett djurs liv .
Något fruktansvärt har hänt .
Hennes ögon blir runda av förvåning .
Tom är en naturlig atlet .
Du säger " dito " , och det är inte detsamma som " Jag älskar dig . "
Tiderna förändras , och vi förändras med dem .
Vi måste tala med dig om Tom .
Vi måste tala med er om Tom .
Vi måste prata med dig om Tom .
Vi måste prata med er om Tom .
Tom har sagt upp sig .
Tom är framåt .
Tom är framfusig .
Tom är artig .
Tom målar .
Tom packar .
Tom ljuger .
Tom är lyckligt lottad .
Tom är för sig själv .
Tom är allena .
Tom är vanvettig .
Tom är vansinnig .
Tom är hungrig .
Tom är hemlös .
Tom är halsstarrig .
Tom är hårdnackad .
Tom är vänlig .
Tom är knäpp .
Tom är hispig .
Tom är stollig .
Tom är färdig .
Tom är lortig .
Tom är smutsig .
Tom är oförskräckt .
Tom är orädd .
Tom är känd .
Tom har rymt .
Tom är förlovad .
Tom äter .
Tom dör .
Tom drömmer .
Tom gråter .
Tom är galen .
Vi är från Ryssland .
Tom lagar mat .
Tom är vid medvetande .
De äter inte kött .
Mamma , var är toalettpappersrullen ?
Någonting fruktansvärt har hänt .
Livet i fängelse är värre än ett djurliv .
Tom är munter .
Tom är glad av sig .
Tom är gladlynt .
Tom fuskar .
Tom är genialisk .
Tom bluffar .
Vad är den turkiska motsvarigheten till meditation ?
Jag har redan sagt det till dig .
Vilket stort hus du har !
Vilket stort hus ni har !
Tom vinner .
Han ser blek ut .
Visa mig var Puerto Rico är på kartan .
Tom behöll min tändare .
Tom gillade den idén .
Tom tyckte om den idén .
Tom bor på en båt .
Tom ser annorlunda ut .
Tom ser äcklad ut .
Tom ser utmattad ut .
Tom ser utpumpad ut .
Tom ser slut ut .
Tom tog ett beslut .
Tom fattade ett beslut .
Tom valde .
Tom gjorde sitt val .
Tom fick mig att göra det .
Tom måste stoppas .
Tom behövde pengar .
Tom behövde kontanter .
Tom kom aldrig tillbaka .
Tom öppnade dörren .
Tom rullade med ögonen .
Tom himlade med ögonen .
Tom satt på trottoarkanten .
Tom blev avvisad .
Tom fick avslag .
Tom fick nej .
Tom fick korgen .
Tom är en sympatisk kille .
Vi måste göra det igen .
Hon är min flickvän .
Vi måste hjälpa Tom .
Vi borde sätta igång .
Vi borde komma igång .
Vi borde ge oss av .
Vi håller kontakt .
Vad har du hört ?
Vad var Toms plan ?
Vad är du bra på ?
När rymde Tom ?
Nu du kommer till Frankrike ska vi åka till Marseille .
Den förra hyresgästen skötte lägenheten utmärkt .
Det är vad alla säger .
Vi värdesätter våra kunder .
Vi klev upp tidigt så att vi kunde se soluppgången .
Vi steg upp tidigt så att vi kunde se soluppgången .
Har du ätit färdigt frukosten än ?
Var är mina saker ?
Var är min golfbag ?
Vem brukade göra detta ?
Vem brukade göra det här ?
Vems idé var det ?
Vems telefon är det där ?
Varför åker inte Tom ?
Varför ger sig Tom inte iväg ?
Skulle Tom gilla det ?
Skulle Tom tycka om det ?
Du kan inte neka det .
Tom var helt hjälplös .
Jag lånade den just .
Jag vet ingenting om hans familj .
Jag vet ingenting om hennes familj .
Jag är i London .
Du är en sådan flörtis .
Njuter du av att förlora ?
Är du rädd för mig ?
Följer du efter mig ?
Följer ni efter mig ?
Kan jag ringa upp dig ?
Kan jag tänka på det ?
Kan jag tänka på saken ?
Har vi råd med det nu ?
Kan du laga en toalett ?
Eld är väldigt farligt .
Jag dricker aldrig öl .
Enligt hans åsikt , ja .
För sent .
Jag kan inte finna min flickväns klitoris .
Behöver ni pengar ?
Var är ni ?
Jag tycker inte om att lära mig oregelbundna verb .
Han var tvungen att lämna skolan för att han var fattig .
Kasta inte bort den här tidningen !
Min farbror bor i New York City .
Tack så mycket .
Vill du äta något ?
Den kalla vinden trakterade luffaren fruktansvärt .
Hans stjärna bleknar .
Målet helgar medlen .
Mitt rum är nummer fem .
Jag vill bara ha kul .
Han ringde mig .
Om jag vore rik , skulle jag åka utomlands .
Jag köpte den igår .
Desto mer man äter , desto mer vill man ha .
Min syster gråter ofta .
Hon rekommenderade kunden en blå slips .
Vilket är ditt favoritnagellack ?
Alla elever i klassen tycker om herr Smith .
Jag är tacksam för din hjälp .
Jag är tacksam för er hjälp .
Skadades någon ?
Gjorde någon sig illa ?
Missade jag någonting ?
Gick det bra i dag ?
Hotade Tom dig ?
Vann du kapplöpningen ?
Vann du kappkörningen ?
Måste jag betala dig ?
Måste jag betala er ?
Har du några kontanter ?
Behöver du någonting ?
Behöver ni någonting ?
Äger du ett handeldvapen ?
Äger du ett eldhandvapen ?
Tom ringer mig nästan varje dag .
Katten är på mattan .
Mittemot stationen .
Han kramade mig .
Vilken tid öppnar marknaden ?
Museet är inte öppet på söndagar .
Dörren stod på glänt .
Tycker du att det är tråkigt här ?
Den filmen var verkligen tråkig .
Jag förstår inte riktigt vad du menar .
Har han accepterat vår inbjudan ?
Jag är fortfarande precis i starten .
Vi upptäckte en hemlig passage .
Har du saknat mig ?
Det är ju en överraskning .
Åh , jag är ledsen !
Mannen som ringde för en timme sedan var Frank .
I byn finns inga tjuvar .
Jag visste inte att hon har ett barn .
Har du tråkigt här ?
Var inte fräck emot mig .
Var inte så dramatisk .
Var inte så negativ .
Var inte så negativa .
Rör inte mina grejor .
Rör inte mina grejer .
Rör inte mina prylar .
Vill du inte åka ?
Rör inte mina saker .
Han berättade aldrig för någon .
Han är rädd för ormar .
Han sjöng vackert .
Hon sjöng vackert .
Hur kan detta vara sant ?
Hur kan det vara sant ?
Hur kan vi tacka er ?
Hur kan vi tacka dig ?
Hur fick Tom reda på det ?
Hur hittade du Tom ?
Hur är detta relevant ?
Hur är det relevant ?
Sjön är stor och vacker .
Det är svårt att sluta röka .
Det är stopp i trafiken på grund av olyckan .
Vilken är starkare , tigern eller lejonet ?
Jag valde mellan två alternativ .
Det var ett extremt grymt krig .
Får jag sitta här ?
Han har på sig glasögon .
Röker du ?
Jag vill inte vila .
Tom är min vän .
Hur lång tid har du på dig ?
Hur lång tid har vi på oss ?
Hur många fick du ?
Hur många fick du tag på ?
Hur mycket vill du ha ?
Hur mycket vill ni ha ?
Jag kan knappt andas .
Jag kan inte sjunga en ren ton .
Jag kan inte komma i kväll .
Jag har varit upptagen .
Det är 99,9 procent effektivt .
Det är nittionio komma nio procent effektivt .
Jag kan inte övertyga Tom .
Jag kan inte heller dansa .
Jag kan inte dansa heller .
Jag kan inte bli inblandad .
Jag hör ingenting .
Jag kan inte höra någonting .
Jag kan inte leva med det .
Jag kan inte riskera någonting .
Jag kan inte ta några risker .
Jag kunde inte bry mig mindre .
Jag skulle inte kunna bry mig mindre .
Jag dödade inte någon .
Jag gör det hela tiden .
Jag tror inte på det .
Jag förtjänar inte detta .
Jag förtjänar inte det här .
Jag har inget emot att hjälpa till .
Jag känner inte igen det .
Jag känner inte igen den .
Jag litar inte på någon .
Jag känner mig väldigt förrådd .
Jag gav inte Tom något val .
Jag fick B i fysik .
Jag fick C i engelska .
Jag antar att du har rätt .
Jag har ryggproblem .
Jag har min egen teori .
Jag har så många idéer .
Jag hoppas att du är hungrig .
Jag behöver bara en minut .
Jag visste att du skulle gilla det .
Jag visste att du skulle gilla den .
Jag visste att du skulle tycka om det .
Jag visste att du skulle tycka om den .
Jag vet allt om dig .
Jag vet allting om dig .
Jag lämnade dig ett meddelande .
När det var mycket kallt , stannade vi hemma .
Jag ser fram emot det .
Jag tappade tidsuppfattningen .
Jag gjorde några ändringar .
Jag tror att Tom ljuger .
Jag tror att vi borde gå .
Jag tror att vi borde åka .
Jag trodde att jag kände dig .
Jag trodde att du åkt .
Jag berättade sanningen för Tom .
Jag förstår helt och hållet .
Du förstår mig .
Vad heter hon nu igen ?
Jag är äntligen färdig med min uppsats .
En snöoväder har dragit in över Sverige .
Nu är vi kvitt .
Jag skulle vilja vara ensam .
Jag skulle vilja hjälpa dig .
Jag skulle vilja följa med dig .
Jag skulle vilja se det .
Jag skulle vilja stå upp .
Jag skulle vilja pröva det här .
Jag är på mitt kontor .
Jag kommer att vara på mitt kontor .
Jag kommer att drömma om dig .
Jag lade märke till att hon satt på främsta raden .
Jag lade märke till att hon satt på första raden .
Vad är lycka ?
" Jag gillar inte morötter . "
" Inte jag heller . "
Ärtor och morötter är vanliga soppingredienser .
Slutligen insåg han sitt misstag .
Patienten var i fara .
Min fru ville adoptera ett barn .
Tror ni att vi kommer att hitta hennes hus ?
Tror du att vi kommer att hitta hennes hus ?
Tom lämnade tv : n på hela natten .
Jag kan inte bara stanna här .
Till slut insåg han sitt misstag .
Jag håller dig informerad .
Jag håller dig à jour .
Jag ringer polisen .
Jag gör mina läxor .
Jag väntar ett samtal .
Jag är glad att du är här .
Jag är så gott som aldrig hemma .
Jag är nästan aldrig hemma .
Jag är här varje kväll .
Jag är här för att hjälpa dig .
Jag är här för att hjälpa er .
Jag kommer inte att dö .
Jag ska inte dö .
Det känns riktigt bra .
Det var ett insidejobb .
Det var ett internt jobb .
Vilken bra tennisspelare Tony är !
Han opererades igår .
I närheten finns ett sjukhus .
Det finns ett sjukhus i närheten .
Jag är .
Det är din tur att diska .
Jag gjorde det igår .
Hur gammal är din farfar ?
Jag var lärare .
Jag tvättade mig .
Giraffer har mycket långa halsar .
Han bad om ett glas vatten .
Vissa fiskar kan ändra sitt kön .
Diplomerade imperialismens lakejer försöker att få en teoretisk grund för sina kannibalistiska praxis i kolonierna .
Förra året bodde jag ihop med David .
Här kommer de .
Titta inte .
Ljug inte .
Hoppa inte !
Fuska inte .
Slåss inte .
Här kommer han .
Hans huvud värkte .
Han går fort .
Det verkar som att han är trött .
Han verkar trött .
Öl är gott .
Tom är svag .
Tom är uppe .
Jag litar på er .
Vissa fiskar kan byta kön .
Den är gjord av läder .
Den är gjord av skinn .
Blunda bara .
Sänk rösten .
Får jag se den där listan .
Låt mig ta en titt .
Mary kom självmant .
Mary kom själv .
Jag har gått och tänkte på det hela dagen .
Jag har tänkt på det hela dagen .
Efter att ha misslyckats två gånger i går vill han inte försöka igen .
John sitter vid Jack .
John sitter bredvid Jack .
Varför ljuger ni ?
Läs inte denna mening .
Din fråga har inget svar .
Er fråga har inget svar .
Spela den sången igen .
Säg åt Mary att jag älskar henne .
Berätta vad du såg .
Talaren är ung .
De närmar sig .
De kommer att ha jättekul .
De är svåra att hitta .
Tom kan inte vara allvarlig .
Tom kan inte vara seriös .
Tom kollade tiden .
Tom kräver uppmärksamhet .
Tom har behov av uppmärksamhet .
Tom dödade inte Mary .
Tom hatar dig inte .
Tom hatar er inte .
Tom hatar inte dig .
Tom hatar inte er .
Tom drack i tystnad .
Tom har dålig hygien .
Tom är miljardär .
Tom är en bra vän .
Tom är neurolog .
Tom är nervspecialist .
Tom är redan där .
Tom är en gammal vän .
Tom är i duschen .
Tom är lång och smal .
Tom tittar på den .
Tom tittar på mig .
Tom är ingen främling .
Tom försvann just .
Tom försvann bara .
Tom försvann precis .
Tom gick just in .
Tom gick precis in .
Tom gick bara in .
Tom vet att han har rätt .
Tom gillar reality-tv .
Tom tycker om reality-tv .
Tom ser frustrerad ut .
Tom gjorde en bra putt .
Tom lovade att hjälpa .
Tom halkade och föll .
Tom låter utmattad .
Tom började skratta .
Tom stal dina pengar .
Tom stal era pengar .
Tom försökte döda mig .
Tom försökte rädda mig .
Tom snavade och föll .
Tom avrättades i elektriska stolen .
Tom gavs en dödande elektrisk stöt .
Tom gick ut och dansade .
Tom kommer att bli överlycklig .
Vi måste göra bättre ifrån oss .
Vi matade just babyn .
Vi matade just barnet .
Vi borde sätta upp en fälla .
Vi är i en konjunktursvacka .
Vi är i en recession .
Vi är i en lågkonjunktur .
Vi är redo för detta .
Hur kan ni inte gilla honom ?
Hur kan ni inte tycka om honom ?
Hur kan du inte gilla honom ?
Hur kan du inte tycka om honom ?
Jag behöver dig .
Tom är ung .
Det är onormalt att äta så mycket .
Ann gillar choklad .
Ann tycker om choklad .
Deadlinen närmar sig .
Här är hon !
Vad har du på dig ?
Vad har du på dig för kläder ?
Vad skriver du ?
Vad för dig hit ?
Vad kan du ge mig ?
Vad kallade du mig ?
Vad kallade ni mig ?
Vad har vi här ?
Vad minns du ?
Vad minns ni ?
Vad mer kan du göra ?
På vintern åkte jag ofta skidor .
Vad mer kan ni göra ?
Exakt vad är det där ?
Vilken årskurs är Tom i ?
Vad var problemet ?
Vad är Toms problem ?
När frågade du Tom ?
Vart är du på väg ?
Var kan jag hitta Tom ?
Vem är redo att beställa ?
Varför sa Tom det ?
Varför sa Tom så ?
Du kan inte ändra på Tom .
Ni kan inte ändra på Tom .
Man kan inte ändra på Tom .
Du kan inte kontrollera mig .
Ni kan inte kontrollera mig .
Man kan inte kontrollera mig .
Du måste göra som jag säger .
Ni måste göra som jag säger .
Talar jag för snabbt ?
Pratar jag för snabbt ?
Är det där mina örhängen ?
Väntar du på Tom ?
Stöter du på mig ?
Är du hungrig över huvud taget ?
Är du fortfarande hemma ?
Är ni fortfarande hemma ?
Luftföroreningar är ett allvarligt globalt problem .
Är du fortfarande gift ?
Är ni fortfarande gifta ?
Kan du inte röra dig fortfarande ?
Skulle jag kunna få en servett ?
Köpte du en nya bil ?
Köpte ni en ny bil ?
Köpte du Tom en hund ?
Köpte ni Tom en hund ?
Köpte du en hund till Tom ?
Köpte ni en hund till Tom ?
Ringde du någonsin Tom ?
Fick du checken ?
Fick ni checken ?
Kände du Tom väl ?
Kände ni Tom väl ?
Tror du på mig nu ?
Tror ni på mig nu ?
Måste du gå nu ?
Måste ni gå nu ?
Måste ni åka nu ?
Måste du åka nu ?
Använder du aftershave ?
Använder ni aftershave ?
Spelar det verkligen någon roll ?
Glöm inte att använda tandtråd .
Droppe blod .
Här är din hund .
Var är min ?
Sådan är lagen .
Han sprang så fort han kunde .
Vem är den där kvinnan i brun jacka ?
Sverige är det största landet i Skandinavien .
Tom såg inte tillbaka .
Det här tåget går mellan Tokyo och Hakata .
En man visade sig i dörren .
Det gör så ont .
Sluta !
Var är min son ?
Tom haltar .
Jag nyser hela tiden .
En man uppenbarade sig i dörren .
Mannen uppenbarade sig i dörren .
Mannen visade sig i dörren .
Glöm inte din väska .
Låt inte Tom se dig .
Låt inte Tom se er .
Se inte så chockad ut .
Tvinga mig inte att göra detta .
Tvinga mig inte att göra det här .
Svara inte på det .
Ödsla inte din tid .
Ödsla inte er tid .
Slösa inte bort er tid .
Slösa inte bort din tid .
Maska inte .
Fyll i den här , tack .
Fyll i denna , tack .
Ta reda på var Tom är .
Var snäll och lämna mig ifred .
Lita inte på honom !
Kanske en annan gång .
Du vet var problemet ligger .
Skulle du kunna lämna mig i fred ?
Amy , du borde gifta dig med honom .
Är perfektion tråkigt ?
Har du rökt ?
Har du sett Tom än ?
Har ni sett Tom än ?
Hur vet du det ?
Hur vet ni det ?
Hur gjorde du det ?
Hur gjorde ni det ?
Hur visste Tom det ?
Hur träffade Tom Mary ?
Hur fick du tag på dem där ?
Hur länge var Tom här ?
Hur många tog du ?
Jag uppskattar hjälpen .
Hon satt och rökte .
Jag ser inget problem med detta .
Han förstod inte hennes skämt .
Jag trodde att vi var bästa vänner .
Häller du upp mer te åt mig ?
Mannen tillstod att det var sant .
Kvinnan beviljades ett stipendium på tusen euro .
Hör och häpna !
Han har dubbelhaka .
Hon har dubbelhaka .
Han sa det med ett flin på läpparna .
Han arbetar inte med något .
Han har inget arbete .
Han har en slapp gångstil .
Hon har en slapp gångstil .
Den där mannen är slapp när det gäller jobbet .
Blomkrukan välte plötsligt omkull .
Vi ses vid femtiden !
Vi ses vid femsnåret !
Parakiten burrade upp sig på pinnen .
Han knäckte nötter .
Hon knäckte nötter .
Spelningen överträffade mina förväntningar flera gånger om .
Han åt en bit av tårtan .
Hon åt en bit av tårtan .
Jag har händelsen i färskt minne .
Friskt vågat är hälften vunnet .
Vi är ingifta släktingar .
Han sprider osanna rykten .
Hon sprider osanna rykten .
Jag klämdes i bilvraket .
I många länder måste man alltid nia främlingar .
Han hade kortklippt hår .
Hon hade kortklippt hår .
Den där kameran tillhör mig .
Bålen syntes långt .
Han rymde långt härifrån .
Han tittade in hos Tom som hastigast .
Hon tittade in hos Tom som hastigast .
Detta är vars och ens ensak .
Jag vill inte ha era hus .
Jag vill inte ha dina hus .
Ingen bryr sig om vad du tycker .
Dina synpunkter är inte av någon vikt alls .
Vem tog hand om hunden medan du var borta ?
Vem tog hand om hunden medan ni var borta ?
Kolet glöd i elden .
Jag älskar min stad .
Välkommen , John !
Vi väntade på dig .
Jag kommer hit varje dag .
Jag kunde inte ljuga för dig .
Jag kunde inte ljuga för er .
Jag bad inte om detta .
Jag bad inte om det här .
Jag flyttade inte på någonting .
Jag sa inget .
Jag sa ingenting .
Jag får inte så mycket post .
Jag behöver ingen hjälp .
Jag konstaterade en sak .
Jag fick reda på någonting .
Jag kom underfund med någonting .
Du gjorde det här med vilje .
Det var söndag i går , inte lördag .
I går var det söndag , inte lördag .
Äter du kött eller är du vegetarian ?
Äter ni kött eller är ni vegetarianer ?
Barnen plaskade glatt i vattnet .
Äntligen börjar molntäcket att lätta .
Han begrep ingenting av det där .
De gick arm i arm i parken .
Jag kikade genom dörrspringan .
Jag knäppte knapparna .
Han talade i vaga ordalag .
Det råder ingen tvivel om det .
Han skrattade sig fördärvad .
Hon skrattade sig fördärvad .
Jag är sprickfärdig av nyfikenhet .
Fågeln vippar på stjärten .
Jag kom inte att tänka på att ta med mig datorn .
Vi fick punktering .
På kvällen var det lite dis i luften .
Han sjöng en sång för att lätta upp stämningen .
Jag får åksjuka .
Jag var tvungen att göra någonting .
Jag fick precis ditt mejl .
Jag fick precis ditt mail .
Jag stötte precis min tå .
Jag stötte precis tån .
Jag visste att jag inte var galen .
Jag visste vad du menade .
Jag visste vad ni menade .
Jag vet hur gammal Tom är .
Jag vet hur detta fungerar .
Jag vet hur det här funkar .
Jag känner Tom personligen .
Jag gillar hur Tom tänker .
Jag tycker om hur Tom tänker .
Jag gillar att vara förberedd .
Jag behöver att du går hem .
Jag gick aldrig och la mig .
Jag gick aldrig och lade mig .
Jag gillar det fortfarande inte .
Jag tycker fortfarande inte om det .
Jag berättar allt för Tom .
Jag tror att Mary tycker om mig .
Jag tror att Mary gillar mig .
Regler är regler .
Vem pratar ?
Jag trodde att jag hörde dig .
Jag trodde att jag var ensam .
Jag trodde att jag var lyckligt .
Jag tyckte att jag var lycklig .
Jag tyckte att det var gott .
Jag tyckte att det var bra .
Jag trodde att du skulle hålla med .
Jag vill tro dig .
Jag vill tro er .
Stäng din bok .
Stäng er bok .
Stäng igen din bok .
Stäng igen er bok .
Skriv aldrig orden " borsjtj " och " sjtji " på tyska !
Jag förstår att Volapük är ett bra språk .
Berings sund avskiljer Asien från Nordamerika .
Jag gjorde det mot min vilja .
Vänligen , mata inte djuren !
Lärare måste förstå barn .
Jag har två utländska vänner .
Jag vågar inte lova någonting .
Inte här !
Jag vet nästan ingenting .
Sluta bete dig som ett barn .
Tom är hemma .
Jag byggde ett hus med utsikt över berget .
Vilka vanor har han ?
Kan du repetera det ?
Man får inte vila på gamla lagrar .
Inte en enda stjärna syntes .
En olycka kommer sällan ensam .
Oaktsamt tal kan få ödesdigra följder .
Mitt bemödande avsatte inget resultat .
Vi är vanliga dödliga .
Vi försökte ta olaterna ur honom .
Tom är sjuk .
Han kom precis i rätt tid .
Han tröttnade på att äta godis .
Han sköt först !
Femtiotvå procent av brittiska kvinnor föredrar choklad framför sex .
En förkylning gjorde honom sängliggande .
Han förbannade sin otur .
Varför beskyller du mig ?
Anklagar du mig för att vara en slöfock ?
Han lindade en filt om valpen .
Kylan ger aldrig med sig här .
Du skulle bara våga röra honom !
Han är ytterst vacker .
Hon är ytterst vacker .
De beviljade medlen förslog inte långt .
Hans skrupelfria agerande gjorde många uppbragta .
Hans svar bestod idel av invektiv .
Hans svar var idel invektiv .
Jag har bott sex månader i Kina .
Han fick ett vederhäftigt svar .
Landet blev till sist oavhängigt .
Han införlivade skämtet med sin repertoar .
Tom använder Windows 7 .
Han har en ganska rustik humor .
Han kände sig föranledd att be om ursäkt .
Han gick i bräschen för att göra byn elförsörjd .
För egen del föredrar jag kaffe framför te .
Själv föredrar jag kaffe framför te .
Tom är sinnessjuk .
Jag pratar arabiska men studerar engelska .
Se upp var du stiger .
Jag kan inte hjälpa dig med det här .
Jag förstår inte vad du säger .
Varför var du frånvarande igår ?
Vad skulle du göra i mitt ställe ?
Se på den där röda byggnaden .
Hur gick du ner så mycket i vikt ?
Jag vill inte dricka nånting kallt .
Vad om han har fel ?
Ser du min bil ?
Var snäll och fortsätt med din historia .
För min del föredrar jag öl framom whisky .
Personligen föredrar jag öl framom whisky .
Jag träffade Mary igår .
De älskar sina barn .
Tom är pensionerad .
Tom har kommit tillbaka .
Jag är trött på att läsa .
Tom skämtar .
Kasta inte nånting på marken .
Samhället består av individer .
Marie följde barnen till skolan .
Varför plågar du mig med det ?
Jag skulle vilja bo i Frankrike .
Det är din tur att sjunga .
Hur gillar ni ert kaffe ?
Jag tror vi är överens .
Tom är mentalsjuk .
Tom är imponerad .
Tom är styvsint .
Jag tror du är svartsjuk .
Han kan varken engelska eller franska .
Har du en reservering ?
Tom är ofarlig .
Tom är oförarglig .
Tom är snål .
Tom sörjer .
Tom är rolig .
Tom är tidig .
Jag vill ha svar och jag vill ha dem nu !
Jag vill ha en förklaring och jag vill ha den nu !
Det är för att du inte vill vara ensam .
Vill du ha nånting att dricka ?
Vill du dansa med mig ?
Tom drunknar .
Jag vill ha en karamell .
Jag vill vara mera självständig .
Tom är i våningen under .
Jag vill se filmen .
Tom är tokig .
Tom är förvirrad .
Tom har erkänt .
Tom är i nedre våningen .
Tom är vid liv .
Tom är på alerten .
Han förklarade den bokstavliga betydelsen av meningen .
Vi lovade .
Vi överlevde .
Vill du ha någonting att dricka ?
Jag tror att vi är överens .
Jag tror att vi håller med varandra .
Jag vill vara mer självständig .
Kasta ingenting på marken .
Personligen föredrar jag öl framför whisky .
För min del föredrar jag öl framför whisky .
Och om han har fel ?
Se upp var du går .
Han verkar snäll .
Jag ska ringa några samtal .
Jag är här för att be om ursäkt .
Jag är bara ärlig .
Jag har sett det här förut .
Jag har sett detta förut .
Det påminde mig om dig .
Det påminde mig om er .
Det är väldigt intressant .
Jane ger aldrig vika .
Jane prutar aldrig på sina anspråk .
Jane ger aldrig med sig .
Lämna min familj ifred .
Håll Tom utanför detta .
Håll Tom utanför det här .
Låt mig ringa min advokat .
Låt mig ta hand om Tom , okej ?
Låt mig tänka en minut .
Låt mig fundera en minut .
Mary är en gold-digger .
Borde inte du gå hem ?
Borde inte ni gå hem ?
Borde inte du åka hem ?
Borde inte ni åka hem ?
Ta ut soporna .
Säg mig vad du tycker .
Berätta för mig vad Tom sa .
Skulle jag kunna få en knäck ?
I år är det jag som har kokat knäcken .
Snön vräker ned utanför fönstret .
Man behöver kramsnö för att göra bra snöbollar .
Det är svårt att bygga snölyktor utan kramsnö .
En lyckad sparktur kräver bra före och ogrusade vägar .
Både is och packad snö är bra underlag för sparkåkning .
Jag har sendrag i benet .
Jag klarade mig helskinnad .
Föreläsningen var verkligen långtråkig .
Han ruskade på huvudet .
Du är så formell .
Jag har ett brokigt förflutet .
Han är ofta borta från skolan .
Han började bli uttråkad .
Hon började bli uttråkad .
Hon är ofta borta från skolan .
Hon ruskade på huvudet .
Jag såg inte en tillstymmelse till ett leende .
Han tyckte att filmen var långrandig .
Hon tyckte att filmen var långrandig .
Hans hobby är styrketräning .
Hennes hobby är styrketräning .
Hans hobby är bodybuilding .
Hennes hobby är bodybuilding .
Bullen var halväten .
Nu är det läggdags för barnen .
Vi är ute med båten .
Bostaden är avlång .
Kursen fortsätter klockan nio .
Hans skjorta är självlysande .
Han tog en uppfriskande promenad .
Hon tog en uppfriskande promenad .
Dessa skor är omaka .
Glaset gick i tusen bitar .
Jag blev genomblöt .
Han har en snusdosa i fickan .
Hon har en snusdosa i fickan .
Han arbetar med att uppteckna traderade berättelser .
Det flitiga bruket av arkaismer tyder på att texten är skriven någon gång under förra seklet .
Jag tycker om te .
Jag kan inte vänta längre .
Han förvirrade oss .
Vad är orsaken ?
Man behöver verkligen inte vara ett stort geni för att översätta från danska till norska ; till och med jag klarar av det .
Att lära sig tala danska är med säkerhet mindre lätt .
Jag har tappat bort min plånbok .
Hela dagen var min pappa på dåligt humör för att han tappat bort sin plånbok .
Denna bok verkar intressant .
Detta är en japansk docka .
Talar du japanska ?
Det var en gång en olycklig , glömsk kille vid namn James , som ständigt förväxlade Mary med Maria .
Därför hatade Maria honom i själ och hjärta .
Att sträva efter sanning är beundransvärt .
Jag vet knappt någonting alls .
Jag vill vinna .
Hon började prata med hunden .
Tom är en desertör .
Tom är en värnpliktsvägrare .
Tom är en helbrägdagörare .
Tom är en urusel dansare .
Tom är på flygplatsen .
Tom är Marys skyddsling .
Tom är Marys protegé .
Han sov tungt .
Han sov djupt .
Hon sov tungt .
Hon sov djupt .
Det finns ingen återvändo .
Det är kallt ute .
Man får aldrig ge upp .
Bara för skojs skull gick jag med på förslaget .
Han spelar golf varje helg .
Det blir för mycket för mig .
Jag behöver sakta ner .
Han var under vatten i tre minuter .
Ge aldrig upp !
Datorn jämförs ofta med människans hjärna .
Det har han inte alls sagt .
Tom är adopterad .
Ett sätt att minska antalet fel i Tatoebas korpus skulle vara att uppmuntra människor att endast översätta till sina modersmål .
Han fick ett raseriutbrott .
Hon fick ett raseriutbrott .
Det är en djupt inrotad tradition .
Han placerade tallrikarna på översta hyllan .
Hon placerade tallrikarna på översta hyllan .
Han är en storätare .
Han är ett matvrak .
Hon är en storätare .
Hon är ett matvrak .
Det närmar sig med stormsteg .
Den närmar sig med stormsteg .
Snoka inte i mina lådor !
Han brast i gråt .
Hon brast i gråt .
Jag är långsynt .
Jag är översynt .
Han hängde sig .
Hon hängde sig .
Han har dålig andedräkt .
Hon har dålig andedräkt .
Regimen störtades till slut .
Han lider av hjärtflimmer .
Han ljög för oss .
Det förklarar varför dörren är öppen .
Hur är det möjligt ?
Du har helt rätt .
Det förklarar varför dörren står öppen .
Han är ful i munnen .
Hon är ful i munnen .
Han var på brottsplatsen .
På bordet står en blomma .
Det står en blomma på bordet .
Hon är tillräckligt gammal för att resa själv .
Han är tillräckligt gammal för att resa själv .
Han är gammal nog för att resa själv .
Tom kan skriva med båda händerna .
Betaler ni tillsammans eller var ock en för sig ?
Vad satsar du på när du lagar mat ?
Förresten såg jag honom igår .
Typisk tjejsnack !
Jag är tacksam över att jag har kunnat koppla av lite .
Han njöt i fulla drag .
Hon njöt i fulla drag .
Nu är det bara att välja mellan allt hon har att bjuda på .
Vad tycker du , vad ska vi hitta på i morgon ?
Jag mår dåligt .
Tack för ditt mejl !
Det vore kul att träffas snart igen .
Hennes tal var för kort .
Tack för mejlet !
Jag mår inte bra .
Du är smartare än vad jag är .
Det doftar gott i huset .
Han brydde sig inte ens om varningarna .
Hon brydde sig inte ens om varningarna .
Jag iddes inte gå dit .
Jag iddes inte åka dit .
Han fick stå i skamvrån .
Hon fick stå i skamvrån .
Kasta inte in handduken .
Han flög upp .
Det var inte en levande själ där .
Det var inte en kotte där .
Han är emot rökning .
Hon är emot rökning .
Han kan inte motstå glass .
Hon kan inte motstå glass .
Känn dig som hemma !
Känn er som hemma !
Han talar alltid emot sig själv .
Hon talar alltid emot sig själv .
Jag är ansvarig för hans beteende .
Han sprang kors och tvärs .
Hon sprang kors och tvärs .
Trädet är grönt .
Tom sänkte rösten .
Tom behöver vinna tid .
Tom lade ned boken .
Tom la ner boken .
Vad sa du till Tom ?
Vad sa ni till Tom ?
Vad berättade du för Tom ?
Vad berättade ni för Tom ?
Vad mer sa Tom ?
Vad mer behöver du ?
Vad händer i morgon ?
Vad är det som pågår här ?
Du behöver bara be om det .
Jag träffar honom ofta .
Håll käften !
Det är ett problem med honom , att han kommer alltid för tidigt .
Låt oss vara ärliga !
Vänta lite !
Stressa inte !
Jag kan inte hålla det för mig själv , hon är verkligen vacker .
Det sägs att han är rik .
Det sägs att han är välbärgad .
Det sägs att hon är välbärgad .
Jag tror knappast det .
Det återstår att se om jag kan komma i tid .
Jag missade att säga att jag inte kan komma .
Inte undra på att presentatören lät konstig , hon var sjuk .
Jag förlorade tålamodet .
Jag tappade tålamodet .
Alltför höga förväntningar är ofta en orsak till besvikelse .
Antingen alla eller ingen .
Allt var förberett i god tid före .
Jag ordnar det .
Han ignorerar mig .
Livet kunde vara en dröm .
Jag bryr mig inte ett skit .
Man vinner ingenting med smicker .
Om du frågar mig , borde vi gå nu .
Flickan stack nyckeln i fickan .
Betalade du för boken ?
Komm tillbaka !
Du bör alltid tänka innan du talar .
När kommer ni att gifta er ?
Berätta det inte för någon !
Jag är ganska nöjd med min nya bil .
Jag har ont i halsen och näsan rinner .
Min fru ringer mig ofta när jag är utomlands .
Jag har inga planer för helgen .
Livet skulle kunna vara en dröm .
Ge mig en torr handduk !
Allting var förberett långt i förväg .
Man bör alltid tänka innan man talar .
Jag kommer med nästa buss .
Vi svängde av åt fel håll .
Såren läker med tiden .
Jag behöver något att skriva med .
I matematik är han ett geni .
Vilken klocka som helst duger , så länge den är billig .
Hjälp !
Hoppa !
Spring !
Stanna !
Vänta !
Vem ?
Vilket skepp var du på ?
Ombord på vilket skepp var du ?
Vad är det som tar så lång tid ?
Vad är det som tar en sådan tid ?
Var har du fått det där ärret ifrån ?
Var kommer det där ärret ifrån ?
Vad gör Tom här ?
Varför gömmer sig Tom ?
Vad är det Tom gömmer sig för ?
När sa Tom det ?
När fick du den här ?
När fick ni den här ?
När sa du det ?
När sa ni det ?
När sa du det där ?
När sa ni det där ?
När behöver Tom den ?
När behöver Tom det ?
Var växte du upp ?
Var växte ni upp ?
Var ska jag lägga den ?
Vems sida är du på ?
På vems sida är du ?
På vems sida är ni ?
Vems sida är ni på ?
Jag kan väl skjutsa dig ?
Varför skjutsar inte jag dig ?
Varför är tåget sent ?
Varför skulle Tom hjälpa oss ?
Man kan inte köpa respekt .
Du kan inte köpa respekt .
Du ser så vacker ut .
Du har slut på ursäkter .
Ni har slut på ursäkter .
Njuter du av det här ?
Njuter du av detta ?
Njuter ni av det här ?
Njuter ni av detta ?
Är du road av det här ?
Är du road av detta ?
Är ni roade av det här ?
Är ni roade av detta ?
Tydligen är jag adopterad .
Kommer ni med oss ?
Kommer du med oss ?
Är du rädd än ?
Är ni rädda än ?
Hotar du mig ?
Hotar ni mig ?
Ring mig när det är färdigt .
Kan någon verifiera det ?
Kan någon intyga det ?
Kan något bekräfta det ?
Kan någon bestyrka det ?
Kan någon bevisa det ?
Kan någon bevisa riktigheten av det ?
Kan jag hämta er någonting ?
Kan jag hämta dig någonting ?
Jag fyller sexton i september .
Jag äter frukost klockan åtta .
Han har ett stort antal böcker .
Hon har ett stort antal böcker .
Jag lämnar böckerna här .
Han föll baklänges .
Hon föll baklänges .
Han föll bakåt .
Hon föll bakåt .
De glömde att låsa dörren .
Hans fru är en synnerligen begåvad kvinna .
Hennes fru är en synnerligen begåvad kvinna .
Det vore bra om du kunde sjunga .
Han studerar dag som natt .
Hon studerar dag som natt .
Kan jag få byta rum ?
Och så levde han lyckligt i alla sina dagar .
Är det bra för hälsan att äta en vitlöksklyfta om dagen ?
Bomull absorberar vatten .
Man måste läsa mellan raderna .
Det var bara en handfull åhörare där .
Vi har i alla fall tak över huvudet .
Han hade hatt på sig .
Hon hade hatt på sig .
Hon stickar avigt .
Han stickar avigt .
Detta är livets skuggsida .
Detta är tröjans avigsida .
Ingen kan förneka detta faktum .
Du är orättvis .
Jag hittade min borttappade plånbok .
Att resa i gott sällskap är alltid kul .
Se ovan !
Jag bor inte i Finland .
De levande kallar jag , de döda begråter jag , åskviggarna bryter jag .
Hen är snygg och smart
Jag vill inte säga hej .
I regel så har män starkare muskler än kvinnor .
Jag pratar med alla er , kompisar .
Jag lär mig i skolan att kvadratroten ur nio är tre .
Har du varit i Mexiko ?
Tokyo är huvudstad i Japan .
Min blodgrupp är A + .
Låt mig hjälpa dig !
Jag behöver inte den här boken .
Jag anlände just .
Hen grät .
Hur många år är du ?
Vad sägs om att gå och simma ?
Det är där borta jag bor .
Skynda dig !
Vi väntar .
Var bodde du nånstans ?
Gillar du snö ?
Tänk på vad jag just sagt dig !
( Åh , vad du måtte känna dig förpliktigad att göra detta )
Jag håller på och äter ett äpple .
Hälsa på Gud !
Wow !
Vad manlig du är !
Du har inte tvättat händerna , inte sant ?
Hur länge stannade du kvar därborta ?
Vi är föräldrar till två barn .
Carla , sångaren , har en magnifik röst .
Jag förstår inte vad du säger ?
Det där är detsamma som hennes hus .
Det var i bergen jag befann mig .
Endast ett språk är aldrig tillräckligt .
Jag började se Namie Amuro .
Ja vad kul , det talas på lojban i Pakistan .
Min pappa bor och arbetar i Tokyo .
Vad slog hen dig med ?
Jag vet att jag är " osvensk " .
Och det tänker jag fortsätta att vara .
Lagom är inte bäst ; bäst är bäst !
Achille föddes 1908 i Paris .
Är det kärlek ?
Mitt yrke är min hobby .
Det lilla kylskåpet är smutsigt .
Tråden är mycket skör .
Jag är inte någon häxa .
Snygg tjej !
Använd den här !
Behöver vi ett universellt språk ?
Hur mycket kostar den dyraste bilen ?
Du ungen , rör inte spegeln !
Tack för att du har förstört min telefon .
Studerar eller jobbar du ?
Småstaden växte och blev till stad .
Det behövs minst tre personer för att leka här .
Jag är en bäbis .
Jag ska hämta upp henne klockan fem .
Det kommer att komma snö .
Jag har ingen cykel .
Hon som jag just nämnde är vacker , betraktad på avstånd .
Hur tog du dig till skolan ?
Hen kan sjunga bra .
Du borde veta .
Var inte orolig , var glad .
Vilka gifter sig ?
Är det så förresten att du spelar fiol ?
Välkommen till mitt hem !
Det här är galet !
Hennes fot upphörde för ett tag att vara henne till nytta .
Jag känner flera elever på den skolan .
Vi borde sticka .
Jag såg honom städa rummet .
Matematik är det ämne jag vill studera sist .
Vilken respektlös typ !
Hon ringde upp mig från Tokyo .
Vad är det här ?
Jag är kroppsarbetande .
Alice är min mamma .
Jag är inte kroppsarbetande .
Jag skulle vilja växla amerikanska dollar till lojbanska rupnu .
Bilen är redo .
Katten gillar att sova bredvid mig .
Det här är min bil .
Det här är inte en mening .
Pojken var tyst .
Hon kunde inte låta bli att skratta .
Skriv ditt namn på listan och ge den till personen bredvid dig .
Jag är alldeles för upptagen för att kunna hjälpa henne .
Pojken höll valpen mot sitt bröst .
Kommer du att stanna hemma en stund inatt ?
Kate och Brian diskuterar målningen .
Är råttan levande eller död ?
Han är född i Schweiz .
Han är schweizisk .
Att veta något om datorer är grunden för alla vetenskaper .
Att tala engelska är inte lätt .
Varför gråter bebisen ?
Jag drömmer mycket .
Vår mamma köpte en hundvalp till oss .
Hon stannade för en stund sedan .
Hon stannade där ett tag .
Hur många äpplen då ?
Språket i ett samhälle är alltid en viktig detalj .
Att vakna är motsatsen till att somna .
Fåglarna flyger .
Du kan prata !
Han är extremt pratsam .
Vad har det med saken att göra ?
Det är värt ansträngningen .
Jag lyckades knappt .
Allt gick fel .
Det är mulet , men det regnar inte .
Jag talar lite spanska .
De där långt där borta är kristna .
Är du buddist ?
Jag förstår inte vad han försöker säga .
Jag förstår inte vad hon försöker säga .
Jag är Alan Tate , Terry Tates son .
Kokade du potatisen med skalet på ?
Hon kom precis i rätt tid .
Detta verk är tidlöst .
Det här verket är tidlöst .
Hans liv saknar mening .
Hennes liv saknar mening .
Han är dum som ett spån .
Hur många gånger om dagen går denna buss ?
Hur många gånger om dagen går den här bussen ?
Han är en man som vi alla respekterar .
Hon erkänner inte att hon har fel .
Han erkänner inte att han har fel .
Hon erkänner sig inte ha fel .
Han erkänner sig inte ha fel .
Kan du passa barnen ?
Hittade de någonting ?
Vet ni vem han var ?
Kan ni passa barnen ?
Gör det dig ledsen ?
Gör det er ledsna ?
Blir ni ledsna av det ?
Få mig inte att döda er .
Ta inga risker .
Slösa inte Toms tid .
Oroa dig inte .
Det är lätt .
Hur mycket kostade den där ?
Jag uppskattar ditt arbete .
Jag uppskattar ert arbete .
Jag kan inte göra det där heller .
Jag kan inte gå till polisen .
Jag kan inte riktigt göra det .
Jag kan inte se någonting .
Jag kunde inte se någonting alls .
Jag fick A på min uppsats .
Jag antar att Tom inte är hemma .
Jag hatar folk som Tom .
Jag hatar människor som Tom .
Jag hatar personer som Tom .
Jag har ett tillkännagivande .
Jag har en kungörelse .
Jag har ett meddelande .
Jag har massor med vänner .
Jag måste göra det själv .
Jag hoppas att det inte är sant .
Jag hoppas att det där inte är sant .
Han ville ha ett bättre jobb än att städa kontorsgolv .
Hon ville ha ett bättre jobb än att städa kontorsgolv .
Jag behöver ett rum för två .
Jag har aldrig ätit kinesisk mat .
Jag har höjdskräck .
Jag skulle gärna ta en kall .
En kall skulle sitta bra .
Den här fågeln finns varken i Japan eller i Kina .
Var vänlig vänta .
Var god vänta .
Efter två minuter tog bensinen i bilen slut .
Efter två minuter fick vår bil slut på bensin .
Andorra är ett litet furstendöme beläget mellan Spanien och Frankrike .
Är du buddhist ?
Hon betedde sig som ett barn .
Vad har hänt med hennes hund ?
Vad har hänt med hans hund ?
Jag byggde ett nytt hus .
Vilken vacker vas !
Jag förstod inte denna fråga .
Jag förstod inte den här frågan .
Jag skulle aldrig tvivla på hans hederlighet .
Jag skulle aldrig tvivla på hennes hederlighet .
Kom på tisdag om du kan .
I dag regnar det .
Det regnar i dag .
Jag beställde denna baddräkt från Frankrike .
Jag beställde den här baddräkten från Frankrike .
Hon spelar golf varje helg .
Varför lyser kattögon i mörkret ?
Varför lyser kattögon i mörker ?
Tom känner inte för att ta med sin hund på promenad den här morgonen .
Tom känner inte för att rasta sin hund den här morgonen .
Hans senaste föreställning var en stor framgång .
Hennes senaste föreställning var en stor framgång .
Han lämnade plötsligt rummet .
Hon lämnade plötsligt rummet .
Följ mig .
Följ med mig .
Följ efter mig .
Det blåste en kall vind .
Min son kom näst sist i mål .
Min son kom i mål näst sist .
Jag kunde bara inte säga nej .
Jag vill bara gå hem .
Jag vill bara åka hem .
Jag vet vad som dödade Tom .
Jag äter bara koscher mat .
Jag borde vila upp mig lite .
Jag borde vila mig lite .
Jag borde få mig lite vila .
Jag trodde att jag förlorat dig ,
Jag trodde att jag förlorat er .
Jag trodde att Tom hade stuckit .
Jag trodde att Tom var död .
Jag trodde Tom var död .
Jag trodde att du gillade mig .
Jag trodde du gillade mig .
Jag trodde att ni gillade mig .
Jag trodde ni gillade mig .
Jag trodde att du tyckte om mig .
Jag trodde du tyckte om mig .
Jag trodde att ni tyckte om mig .
Jag trodde ni tyckte om mig .
Jag trodde att du var Tom .
Jag är bara en taxichaufför .
Jag har varit där mycket .
Det är nästan omöjligt .
Det är närapå omöjligt .
Kom ned från scenen bara .
Tom kommer inte överens med sina grannar .
Bort med tassarna !
Håll dina händer borta från mig .
Han knäckte ryggen på boken .
Kinesiska tidningar övervakas av regeringen som behåller rätten att ändra innehåll för att passa den rådande partilinjen .
Hon spelar Monopol .
En skola i Storbritannien har frångått läroböcker till förmån för iPads i klassrummet .
Sluta vara så dramatisk .
Jag misstog mig .
Jag tog fel .
Jag vet att pengar inte är allt .
Han gör allt som står i hans makt .
Hon gör allt som står i hennes makt .
De tog skada för livet .
De fick men för livet .
En sten föll från hans hjärta .
En sten föll från hennes hjärta .
Vår galax heter Vintergatan .
Talar ni bulgariska ?
Hon har något emot rödhåriga .
Jag såg henne städa ett rum .
Denna förordning träder i kraft från och med nästa år .
Alla goda ting är tre .
Du gissade rätt .
Boken var fortfarande i bilen .
Mitt löfte att komma nästa måndag håller fortfarande .
Det finns vissa nackdelar .
Koppen är på bordet .
Jag älskar den här koppen .
Kartan hänger på väggen .
Det här är min fru , Minna .
Han läser en bok .
Säg att du skämtar !
Katten satt på mattan .
Tom kunde inte hitta Mary .
Tom kunde inte finna Mary .
Tom fritog gisslan .
Tom har inget perspektiv .
Tom håller i en kniv .
Tom är på sjukhuset .
Tom är bara rädd .
Tom är på väg hit .
Tom är fortfarande skeptisk .
Tom har någonting på gång .
Tom väntar på dig .
Tom väntar på er .
Tom lever ett stillsamt liv .
Tom lånade mig den där DVD : n .
Tom hade aldrig en chans .
Tom hade aldrig någon chans .
Tom sköt mig i benet .
Han kom till Japan för sju år sedan .
Batterierna i min miniräknare är slut .
Hon är ungefär lika gammal som jag .
Jag tycker om sashimi .
Vad bra han spelade !
Han skriver till mig varje vecka .
Jag ångrar inte vad jag har gjort .
Jag ångrar inte det jag gjorde .
Är de amerikaner ?
" Hur mycket är klockan ? "
" Hon är halv elva . "
Han pratade bara dumheter .
Detta är inget att skratta åt .
Hon körde in bilen i garaget .
Jag ser ut som en ren .
Jag lovar , det är värt ansträngningen .
Jag kan inte vara lugn .
På stranden kan man tillbringa tid med sina vänner .
Toms förklaring är mycket detaljerad .
För vem ringer klockorna ?
Hon hade en röd baddräkt på sig .
Skulle du vilja ha ett kokt ägg till frukost ?
Gamla vänner kontaktade mig .
Du bör låta din son bli självständig .
Trafikhinder varade i en timme .
Trafikstockningen varade i en timme .
Om det är gratis , ta så mycket du kan .
Denna bok innehåller många vackra bilder .
Öppna inte dörren innan tåget har stannat .
Ditt hår är för långt .
Han har en hel del kreativa idéer .
Taket på huset läcker .
Han var tvungen att lämna skolan för att han var medellös .
Släng inte den här tidningen !
Jag tror inte att de accepterar dessa villkor .
Han kommer snart .
Jag slutade röka för ett år sedan .
Jag vill skicka det här brevet till Japan .
Bara ät , om du är hungrig !
Koppen står på bordet .
Där är en pojke .
Pojken har en tidning .
Vi bor i Puistokatu .
Också detta är ett äpple .
Han ville absolut börja gräla .
Järn leder värme bra nog .
Tala tydligt !
Jag hade pluggat engelska i två timmar när han kom in .
Jag tycker det är bäst att vi skippar cyklingen .
Han misstänktes vara spion .
De erbjöd assistans .
De erbjöd hjälp .
Fotboll är populärare än tennis .
I dag ska jag gå på konsert .
Jag skulle vilja se den .
Om jag vore du så skulle jag inte bry mig om det .
Det här teet smakar gott .
Jag har väntat i nästan en halvtimme .
Vi motsätter oss krig .
Vi är emot krig .
Har du någonsin varit utomlands ?
Är ni ägaren av detta hus ?
Är ni detta hus ägare ?
Är ni det här husets ägare ?
Vad svarade du ?
Annars måste vi annullera den här beställningen .
Han kan tala franska och engelska .
Han var väldigt trött .
Himlen är oskyldigt blå .
Jag är ursinnig .
Jag är rasande .
Hunden är smart .
Jag älskar äpplen .
Jag gillar att simma .
Jag tycker om att simma .
Jag tycker om simning .
Jag tycker om tennis .
Jag har en vän i England .
Jag har en kompis i England .
Jag är säker på att han kommer .
Jag är säker på att hon kommer .
Kan du ens föreställa dig hur mitt liv är ?
Kan du ens föreställa dig hurdant mitt liv är ?
Vad sa mannen ?
Två plus två är fyra .
Du skulle inte ha behövt ta taxi .
Bröder !
Han rördes till tårar .
Hon rördes till tårar .
Ge mig ett glas mjölk .
Jag tycker inte om dig längre .
Hunden heter Ken .
Han kan ha gått en annan väg hem .
Jag tycker om äpplen .
Jag gillar äpplen .
Han är stolt över att vara doktor .
Han är stolt över att vara läkare .
Dagen randas .
I esperanto slutar alla substantiv på o .
Vad lagar du ?
Han hittade min cykel .
Jag måste stryka min skjorta .
Min storebror är lärare .
Jag lyssnar på Björks senaste låt .
Vi skulle vilja ha en flaska rosé .
Jag har glömt min PIN-kod .
Jag vill inte översätta den här meningen .
Jag vill inte översätta denna mening .
Byggdes denna mur för att hålla människor ute eller för att hålla dem inne ?
Byggdes denna mur för att hålla människor ute eller inne ?
Byggdes den här muren för att hålla folk ute eller för att hålla dem inne ?
Jag svimmade .
En polygon har många vinklar och lika många sidor .
Alt övrigt kolla upp i Wikipedia !
Jag skulle göra vad som helst för kärlek .
Jag skulle göra vad som helst för kärleken .
Det är bara en droppe i havet .
Det är inte något allvarligt .
Ditt rum är väldigt stort .
Ditt hus är stort .
Ert hus är stort .
Ormar äcklar Lisa .
Jag bor på Malta .
Rökning är strängt förbjudet här .
Sätt dig ned och känn dig som hemma !
... sa flickan !
Det är svårt att tala offentligt .
Om han är utomlands , har han ständigt hemlängtan .
Han ville smickra mig .
Hon ville smickra mig .
Blir du nervös om du måste tala inför många människor ?
Jag är fri som en fågel .
Det var en stor förlust för mig .
Det kan vara sant .
Det finns inte ett enda moln på himlen .
Jag skyller på ditt skägg .
Han bor inuti ett äpple .
Ett språk är en dialekt med en armé och en flotta .
Han längtar ständigt hem när han är utomlands .
Hon längtar ständigt hem när hon är utomlands .
Jag har ett par med päron .
Nu ska du få höra min hemlighet .
Den är mycket enkel : Det är bara med hjärtat som man kan se ordentligt .
Det viktigaste är osynligt för ögonen .
Hur tar jag mig dit bäst ?
Han kommer tillbaka sex .
Du sa att du var lycklig .
Ni sa att ni var lyckliga .
Tom åt någonting .
Jag vill bara veta .
Klava överförenklar allting .
De är ivriga på att få veta vad som hände .
De är spända på att få veta vad som hände .
Det är ett extremfall .
Vi har large , medium och small .
Vilken storlek vill du ha ?
Vi har large , medium och small .
Vilken storlek vill ni ha ?
Tom tog av sig skjortan .
Tom tog av sig tröjan .
Tom försökte behålla lugnet .
Tom ville träffa Mary .
Tom är för tidigt född .
Du stötte på honom tidigare , eller hur ?
Ni stötte på honom tidigare , eller hur ?
Vill ni spela tennis med oss ?
Vill du spela tennis med oss ?
Enligt lag har Liisa rätt till skadestånd .
Tom kunde inte kontrollera sig själv .
Nu är goda råd dyra .
Han tvärstannade .
Hon tvärstannade .
Han tvärbromsade .
Hon tvärbromsade .
Han tvärnitade .
Hon tvärnitade .
Den här sjön är verkligen fiskrik .
Den här sjön är verkligen rik på fisk .
Han har en skruv lös .
Hon har en skruv lös .
Du måste hjälpa henne .
Ni måste hjälpa henne .
Jag såg på honom att han bara låtsades läsa .
Han tog med sig en kompis .
Han tog med sig en vän .
Mitt språk är inte med på listan !
Jag måste springa ärenden .
Klandra inte mig !
Jag har inte något att göra med den där videon .
Festen var så tråkig att jag tog till flykten nästan omedelbart .
Att sträva mot strömmen kräver mod .
Det var allt annat än trevligt .
Det finns all anledning att betvivla att det är sant .
Jag försökte att undanröja alla tvivel .
På era platser , färdiga , gå !
Jag beklagar att jag inte gick dit .
Detta är mycket typiskt för dig .
Det kan ingen motstå .
Det är inget att klaga på .
Tack för skjutsen .
Det kan du lita på .
Får jag besvära Er med en anhållan ?
Han fyllde glaset med vin .
Vad behöver du veta ?
Vad måste du veta ?
Han spetsade öronen .
Hon spetsade öronen .
Han hade öronen på helspänn .
Hon hade öronen på helspänn .
Han är den självgodaste människa jag känner .
Hon är den självgodaste människa jag känner .
En tår tillrade ned för hans kind .
Jag ångrar att jag inte åkte dit .
Jag ångrar att jag inte gick dit .
Skyll inte på mig .
Jag har ingenting att göra med den där videon .
Min bil är tysk .
Åh herregud !
Vem arbetar ikväll ?
Var nu inte så skadeglad !
Det var en bra idé .
Gör det aldrig igen !
Kan du simma alls ?
Låt inte folk göra dig galen över pengar , hår och kläder .
Varje fredagskväll gick de och drack sig fulla .
Jag minska mängden ätit godis .
Jag minskar på godisätandet .
Var är dina nycklar ?
Han gör ingenting annat än klagar dagarna i ända .
Skulle du vilja ha ett glas vatten ?
Är din fru kvar i Amerika ?
Är din fru fortfarande i Amerika ?
Det är värt ett försök .
Han tycker inte om kaffe .
Brott lönar sig inte i längden .
Kriminalitet lönar sig inte i längden .
Kriminalitet lönar sig inte i det långa loppet .
Kriminalitet lönar sig inte på lång sikt .
Jag var försenad på grund av trafiken .
Vilken bra idé !
Vi hörs .
Jag skulle gärna vilja ha en bit ost , tack .
Hon litade på mig .
Hon kan inte bara prata engelska utan också franska .
Hon kan inte bara tala engelska , utan också franska .
Jag äter ett äpple .
Ursäkta , var ligger posten ?
Alla i Tyskland har rätt att vistas ute i naturen .
Ni vet att vi inte har så mycket tid just nu .
Hela den polska östersjökusten utgörs av sandstränder .
Hon tycker inte om sport och det gör inte jag heller .
Hon tycker om vin .
Hon gillar vin .
Jag går sällan på bio .
Jag tror killen menar allvar .
Oj , vad synd .
Var och en kan naturligtvis ha en annan åsikt .
Glöm det , det blir inget !
Det kan man tycka annorlunda om .
Jag tror att den här killen menar allvar .
Tom vill inte bli läkare , trots att han är väldigt på naturvetenskap .
När såg du henne senast ?
Tom skrattade åt alla Marys skämt .
President Truman var tvungen att fatta ett svårt beslut .
President Truman var tvungen att ta ett svårt beslut .
Tom har dörrarna låsta om natten .
Fler och fler studenter ansluter sig till protesterna .
Jag undrade bara om du har lyckats hitta någonstans att bo .
En av dina knappar har lossnat .
Till följd av konstant hunger och utmattning dog hunden till slut .
Men när jag försökte vrida duschkranen rann en svart , bubblig vätska ut .
Varorna som beställdes från England förra månaden har inte anlänt än .
Laurie älskar mig .
Hur fick du tag på en sådan stor summa pengar ?
Skynda dig tillbaka .
Varför skulle Tom vilja hjälpa oss ?
Låt oss sköta vårt jobb .
Tom kan inte bestämma sig för vad han ska köpa .
Han fick sitt vänstra ben skadat i en olycka .
Orsaken till olyckan är okänd .
Regnet slog emot fönstren .
Han var riktigt kall .
Vi har saker att göra .
Han kan inte ha tappat bort sina nycklar .
Han är världens rikaste man .
Han skulle aldrig få se sina föräldrar igen .
Det var väldigt svårt .
Jag är redan sen .
Jag äger två böcker .
Var är hon ?
Det är inte alltid lätt att skilja på japaner och kineser .
Telefonen är trasig .
Experimentet var lyckat .
När ska du åka till Europa ?
Han har ingen biljett .
Hon har ingen biljett .
Han är lagkapten .
Tala högre så att alla kan höra dig .
De är lika starka som vi .
Tåget är försenat på grund av snön .
Tåget försenades av snön .
Du tycker verkligen om att äta .
Du gillar verkligen att äta .
Så hur gick det ?
Blev det någon fisk ?
Kan du se dem ?
Kan ni se dem ?
Jag tappade lusten .
Han har tappat lusten .
Han har ingen lust att gå på bio .
Han har ingen lust längre .
Det finns ingen anledning till all denna uppståndelse .
Hur kommer det sig att du har tappat lusten ?
Hur kommer det sig att du inte har någon lust längre ?
Hon hade ingen lust att följa med till affären , så hon stannade hemma istället .
Har du lust att följa med i morgon ?
Jag har lust att gå på bio i morgon .
Jag skulle gärna följa med dig och shoppa , men jag har läxor att göra .
Spärra utgångarna !
En snövall blockerade utfarten .
Ingenting kan hindra oss nu .
Källaren är översvämmad .
Den här bäcken svämmar över varje vår .
Han gick planlöst omkring på stadens gator .
Passa på att njuta av stillheten .
Skulle vi kunna få lite tystnad här ?
Vi har varit strömlösa i tre dagar nu .
I morgon kommer vi att ha varit strömlösa i tre dagar .
Han glömmer aldrig att betala en räkning .
Han ådrog sig en tillrättavisning .
Halva deras årsinkomst går till mat .
Plankorna var delvis täckta av en presenning .
Lämna dörren på glänt när du går .
Han tycker om löskokta ägg .
Han gillar löskokta ägg .
Hon stiger ofta upp mitt i natten för att äta .
Hon kliver ofta upp mitt i natten för att äta .
Han låtsades hålla med henne .
Allt var bara tomma ord .
Han låtsades hålla med om att det var en bra plan .
De har inte acklimatiserat sig än .
De är fortfarande ovana vid klimatet .
Du ska ta tre tabletter fem gånger om dagen .
Du ska ta tre tabletter fem gånger dagligen .
En stor isklump for ned från taket och träffade marken med en hög duns .
Det är bara ett insektsbett .
Han tröttnar aldrig på att äta godis .
Ser jag verkligen så sorgsen ut ?
Vi måste utarbeta en plan .
Den här filmen är väldigt svår att få tag på just nu .
Man planerar att uppföra ett kraftverk precis här .
Han måste vara någonstans i pensionsåldern .
Hon har ett tjockt lager smink på sig .
Desto längre söderut man kommer , desto mildare blir klimatet .
Hon studerar filosofi på landets förnämsta universitet .
Skulle jag kunna få låna om den här boken ?
Går det att låna om den här boken ?
Går det att förlänga lånetiden på den här boken ?
Ingenting är säkert när det gäller honom .
Är dessa däck slirfria ?
Dubbdäck är förbjudna på den här gatan .
Utan dubbdäck tar du dig inte upp för den där backen .
Vi har inte hela dagen på oss .
Det är lugnt .
Sätt dig ned och andas en stund nu .
Jag har inte en muskel på hela kroppen .
Han är muskulös .
Kan vi inte bara spankulera runt i parken ?
De flanerade en hel eftermiddag på stan .
Jag luras aldrig .
Han blev förd bakom ljuset .
Flickan är nu utom fara .
Patientens skador är inte livshotande .
Patienten har inga livshotande skador .
Patienten vårdas på intensiven .
Han täljde en grillpinne med sin fickkniv .
Man får ta vad man har .
Hon är gammal och erfaren .
Är du helt säker på din sak ?
Jag får väl gå och ta reda på det själv .
Det är ett helt outforskat område .
Han har ett gott hjärta .
Hon har ett gott hjärta .
Han gjorde det helt på eget bevåg .
Jag kan inte minnas hans namn .
Jag kan inte komma på hans namn .
Jag kommer inte på hans namn .
Jag minns inte vad han heter .
Jag kan inte minnas vad han heter .
Jag kan inte komma på vad han heter .
Jag kommer inte på vad han heter .
Jag är ekonomiskt självständig från mina föräldrar .
Jag har hört att de har god service på den här restaurangen .
Partiet påstår sig tjäna folket .
Är den här burken helt tätförslutande ?
Säg inte att du har glömt passet hemma .
Min katt älskar räkor .
Den här terminen har hon gjort ytterligare framsteg .
Nu slog vi två flugor i en smäll .
Hackar du grönsaker ?
Tiden är ännu inte mogen .
Han vet alltid vad som är på modet .
Hunden åt upp sin mat och slickade sig om nosen .
De ska lansera en ny produkt nästa vecka .
Visa vad du går för !
Vi ska gå på en förhandsvisning nästa vecka .
I dag förhandsvisar vi " The Hobbit " i stora salongen .
Han spände ut bröstkorgen .
Han skummade igenom texten .
Jag är hungrig som en varg .
De tände en myggspiral .
Sådana här starka laserpekare är förbjudna på allmän plats .
Förlåt , det hade jag fullständigt glömt bort .
Skillnaden är i en princip obefintlig .
Det kommer fler tillfällen , jag lovar .
Det gör lite ont precis här .
Men det är ju absurt .
Varför säger du inte det här förrän nu ?
Värmeljusåtgången hemma hos oss är galet hög .
Det går åt galet mycket värmeljus hemma hos oss .
Skulle du kunna hålla en plats åt mig ?
Om du inte vet svaret , försök att chansa .
Stäng fönstret , så att du inte blir förkyld .
Han har gått ur tiden .
Det var ett känslofyllt möte .
Nu hade du flax .
Nu hade du allt bra tur .
Jag kommer att sakna dig .
Du är saknad här hemma .
Han har en självlysande pyjamas .
När jag var liten hade jag en självlysande pyjamas med skelett på .
Hajar du ?
Han fattade ingenting .
Hur skulle definiera det här ordet ?
Han stod vid dörren .
De offentliggör resultatet i morgon eftermiddag .
Säg inte ett knyst .
Han sa inte ett knyst .
Enstaviga ord är lätta att komma ihåg .
Enstaviga ord är lätta att blanda ihop .
På plats var en handfull åhörare .
Han blev mobbad i skolan .
Hon trängde sig fram i folkmassan .
Skrivbordsarbete är ofta monotont .
Nu är det färdigdukat .
Ser du till att bordet är färdigdukat när gästerna kommer ?
Han sitter vid datorn .
Två demonstrationer hölls på torget i helgen .
Hur lång garanti är det på datorn ?
Först måste vi skrapa bilrutorna .
Han skrapade bilrutorna .
Nu har hela bilen immat igen .
De har köpt nya högtalare .
Hur mycket kostade ert högtalarsystem ?
Från honom får man alltid bara undvikande svar .
Med denna inspelning kan vi få dem att göra vad vi vill .
Björnen brummar .
Jag får alltid ont i axeln när jag springer .
Vi har bara en stump kvar .
Han läste boken i ett streck .
Självgodare människa får man söka efter .
En mer egoistisk människa får man söka efter .
En dyrare restaurang får man söka efter .
Nu får du ta och skärpa dig .
Hur ofta kollar du din mejl ?
Pesto är Guds gåva till folket .
Han är en god människa .
Jag har inte ätit soppan och jag kommer inte att göra det .
Jag är ledsen att jag har inte skrivit till dig på så länge .
Den här cd kostar tio dollar .
Tom har två söner .
Båda av dem bor i Boston .
Titta på huset med det röda taket .
Tom har två sönder .
Bägge bor i Boston .
Abborren är vanlig i svenska insjöar .
Hon kände sig föranledd att abdikera .
Vad har du för telefonabonnemang ?
Hur stor del av fakturan består av abonnemangsavgift ?
Antalet abonnenter har fördubblats de senaste fem åren .
Vi har abonnerat en buss .
Bussen är abonnerad .
Hon har precis genomgått en abort .
Abortfrågan är stor just nu .
Sveriges abortlagar är inte särskilt restriktiva i jämförelse med andra länders .
Han är absolutist .
Vår filosofi vilar på absolutistiska grunder .
Trasan absorberade vätskan .
Han har abstinens .
Har du skrivit färdigt ditt abstract än ?
De sjunger a cappella .
Efter stoppet accelererade tåget snabbt .
Var ligger accenten ?
Han kan inte skilja på ett accenttecken och en apostrof .
Detta är inte acceptabelt .
Han kommer inte att acceptera denna behandling länge till .
Utan accessoarer känner jag mig naken .
Piano och gitarr är vanliga ackompanjemangsinstrument .
Kören ackompanjeras av Emil på piano .
Alla anställda jobbar på ackord .
Han har ackordlön .
De tittade på en actionfilm .
Vilken är din favoritactionrulle ?
Han klarar inte av addition , än mindre multiplikation .
Vi måste komma på en ad hoc-lösning .
Han är adlad .
Hur hög är administrationsavgiften ?
De adopterade två barn från Asien .
Han arbetar på en adoptionsbyrå .
Vad har du för adress ?
Paketets adressat har fortfarande inte hämtat ut sitt paket .
I fönstren lyser adventsljusstakarna .
Hon hängde upp en röd adventsstjärna i fönstret .
Vet du vad årets adventskalender är ?
Jag är arg .
Det sista tåget har redan farit .
Det sista tåget har redan åkt .
Ni är orättvisa .
Lägg inte plånboken ovanpå elementet .
" Aeroplan " är ett nu föråldrat svenskt ord för flygplan .
Han har drabbats av afasi .
Han drabbades tidigt av afasi .
Skoterns affektionsvärde överstiger dess pengavärde .
På denna vägg är affischering förbjuden .
Hon äger en trevligt liten affär i Gamla stan .
Han arbetar som affärsbiträde .
Han blev påkommen med att avslöja affärshemligheter .
Tror du på min affärsidé ?
Hon har kommit på århundradets affärsidé .
Han studerar affärsjuridik .
Han gjorde en Afrikaresa tidigt förra våren .
Han använder alltid en exklusiv aftershave .
Han använder alltid en exklusiv after shave .
Ska ni med på afterski i kväll ?
Ska ni med på after ski i kväll ?
Glöm inte att det är afterwork i kväll .
Glöm inte att det är after work i kväll .
Barnaga är förbjudet i Sverige .
Barnaga är fortfarande tillåtet i många länder .
Vad står på dagens agenda ?
Vi måste agera nu .
Det finns ingen anledning att hysa agg emot honom .
Hon är aggressiv .
Hennes hund går på agility .
Han är agnostiker .
Han lider av agorafobi .
Partiet lämnade agrarpolitiken bakom sig för länge sedan .
Det kom som en aha-upplevelse .
För henne var det en aha-upplevelse .
Är bilen utrustad med airbag ?
Ajabaja !
Den rör du inte !
Genom att läsa nättidningen håller sig morfar ajour .
Han är akademiledamot .
Han lever på a-kassa .
Alla har en akilleshäl .
IKEA är en akronym för Ingvar Kamprad Elmtaryd Agunnaryd .
Akta dig för henne !
De ska sälja sina gamla möbler på aktion .
De ska aktionera ut sina gamla möbler .
Har du aktiverat virusskyddet ?
Virusskyddet är aktiverat .
Alla barn behöver aktiveras .
Denna fråga är ytterst aktuell .
Han arbetar som akupunktör .
Hur akut är det ?
Han fick åka in på akuten .
Detta är ett akutfall .
Väl inne på akutmottagningen sa de att han bara hade inbillat sig allting .
Den här mannen behöver akutvård .
Hon målar med akvarellfärger .
En vecka senare inflöt en alarmerande rapport .
Det här blir hennes tredje album .
Trots att han är nittio år är han fortfarande mycket pigg och alert .
Det gäller att vara på alerten om man inte ska missa någonting .
Hon lider av alexi .
Har han alibi ?
Alkemi är en utdöd vetenskap .
Han har lovat att han ska ta tag i sitt alkoholberoende .
Är den här drinken alkoholfri ?
Har ni något alkoholfritt ?
Hon har sagt upp bekantskapen med sin alkoholiserade mamma .
Denna bil är försedd med alkohollås .
Den här bilen är utrustad med alkolås .
Han har dåliga alkoholvanor .
Lägenheten har en alkov .
Allemansrätten tas för givet av många svenskar .
Har du ingenting att säga ?
Har du inte någonting att säga ?
Vi måste köpa en ny router .
Jag är längst i vår klass .
Hans sjukdom orsakas av överdriven alkoholkonsumtion .
Köpenhamn är Danmarks huvudstad .
Jag beundrar verkligen ditt mod .
Om du tror att det var mitt fel är du inne på fel spår .
Resultatet var värt noll .
Det var kul att höra .
Detta kan inte beskrivas med ord .
Ditt förslag låter bra .
Köpenhamn är huvudstaden i Danmark .
Du var min räddare i nöden .
Om ditt sinne matar ditt svärd , kommer ditt svärd säkerligen att äta ditt sinne .
Erfarenheten räknas .
Erfarenheten har visat : pengar ger inte lycka .
Erfarenhet lönar sig .
Hur kunde jag trösta dig ?
Hon glömde att mata hunden .
Hon hade goda skäl att söka skilsmässa .
Du behöver bara be om den .
Vår son dog i kriget .
Tom drack en hel del vodka under sin resa till Ryssland .
Kan jag äta denna kaka ?
Du måste hålla dig i form .
Stoppa tjuven !
I detta avseende , har du rätt .
Sluta skratta !
Det låter bra !
Saken stör mig fortfarande .
Jag tycker att det är fantastiskt .
Jag hoppas att alla dina drömmar blir verklighet .
Vid midnatt skall jag gå fram genom Egypten , och allt förstfött i Egyptens land skall dö .
Ju förr desto bättre !
Därefter var jag alldeles slut .
Det lönar sig nog att vänta .
De håller på att äta just nu .
Han är en bra talare .
Egentligen ville Liisa gå ut och festa , men hon stannade hemma .
Egentligen får man inte vänsterprassla .
Hörde ni mig inte ?
Vi använder endast tio procent av vår hjärna .
Vi kan inte låta Tom dö .
Det finns ingen gratis lunch .
Du klarade det !
Jag vet att det inte är lätt .
Han är mycket oförskämd .
Hans ansikte strålade av lycka .
Hur gammal är din farbror ?
Detta bolag har hittills varit synnerligen framgångsrikt .
Killen är oförskämd .
Detta är långt ifrån säkert .
Det var inte det jag letade efter .
Det är självklart .
Från månen , kunskap .
Från stjärnorna , kunskap .
Den där typen vet inte hur man beter sig .
Han är väldigt oförskämd .
Hur gammal är din morbror ?
Du lyckades !
Du gjorde det !
Han är din vän .
Han är din kompis .
Han är din kamrat .
Jag tror att det skulle vara roligare att gå tillsammans .
Han blev väldigt rädd .
Under kvällen kommer det att sluta snöa .
Han menar det på allvar .
Muntra upp dig !
Kosta vad det vill !
Kort och gott .
Kosta vad det kosta vill .
Liisa anklagade mig för vårdslöshet .
Ryck upp dig !
Ryck upp er !
Vill du ha en snigel på ögat ?
Var är den grekiska ambassaden ?
Han har två bilar .
Hon talar portugisiska .
Hon vill ha någonting väldigt speciellt på födelsedagen .
Jag är förvånad att han antog erbjudandet .
Jag är förvånad att han accepterade erbjudandet .
I morgon kommer jag inte att vara här .
I morgon är jag inte här .
Damaskus ligger i Syrien .
En sten föll från mitt hjärta .
Tack för lånet .
Vem är din lärare ?
Du måste absolut följa med !
Slå upp numret i telefonboken !
Ta inte illa up !
Ingen orsak !
Det är bara att ta !
Parkering förbjuden !
Sköt om dig !
Har du ett problem , är det ibland bättre att vara praktisk och sättä igång med lösningen än att fundera ändlöst .
Hämnden är ljuv .
Prata inte dumheter !
Han är inne .
Han sa ja .
Vädret är sämre i dag än i går .
Han sade ja .
Prata inte smörja !
Sätt igång !
Liisa jobbar och studerar samtidigt .
Inga skämt , tack !
Det går upp för mig .
Man får inte bryta sitt löfte .
Liisa är benägen att gråta på bio .
Lägg dig inte i det här !
Försök inte att undvika ansvar !
En empatisk flicka kan känna med en väns känslor .
Under tiden kan jag göra mig förstådd .
Somalia heter " as-Sumal " på arabiska .
Glöm det !
Var inte så hård mot dig själv !
De roade sig med video-spel .
Du måste förbereda dig för det värsta !
I matematik var han vida överlägsen alla andra .
De roade sig med att spela tv-spel .
Försökt inte att fly från ansvar .
Liisa studerade vid sidan av jobbet .
Vad är du rädd för ?
Vad är ni rädda för ?
Vad har vi för val ?
Vad tycker du , Tom ?
Vad är alternativet ?
Vad heter Tom i efternamn ?
Vad är det för fel med det ?
Vad hette du nu igen ?
Vad var det du heter nu igen ?
Var är bilnycklarna ?
Var är Toms saker ?
Var kom den ifrån ?
Var kom det ifrån ?
Var hittade du Tom ?
Var fann du Tom ?
Var fick du tag på den där ?
Är du fortfarande arg på mig ?
Är ni fortfarande arga på mig ?
Var trevligare mot din syster .
Var trevligare mot er syster .
Sa någon någonting ?
Såg du den på riktigt ?
Såg du det på riktigt ?
Hittade du din handväska ?
Hittade du din börs ?
Min vän är sjutton år .
Min kompis är sjutton år .
Kan vi inte spela tv-spel i kväll ?
Bär hit bordet .
Ta tag i varsin ände och bär hit bordet .
Ni behöver inta vara rädda .
De håller ihop som klister .
Tom undrade om det som Mary sade var sant .
Hon var en riktig pärla .
Är ditt modersmål kinesiska ?
Är kinesiska ditt modersmål ?
Något sådant kan hända vem som helst .
Sådant händer ju ibland .
Jag sätter mig så länge .
Sådant händer .
Koncentrera dig på ditt uppdrag !
Koncentrera dig på vårt uppdrag !
Absolut förbjudet .
För att vinna tid tog vi planet .
Jag vill inte orsaka några olägenheter .
Är detta äkta silver ?
Var uppriktig mot mig .
Det var ett till synes genuint leende .
Det knackade på dörren .
Det knackar på dörren .
Dörrklockan ringde .
Någon ringde på dörrklockan .
Det är hans omedgörlighet som irriterar mig .
Mormor har gjort en rulltårta .
Vi vill rösta .
Det börjar bli dags att börja .
Det är ingen brådska .
Hajar är goda simmare .
Behöver du dricka vin ?
Varför har koalor ingen navel ?
Föredrar du en manlig eller kvinnlig doktor ?
Jag tar det .
Mina ögon gör ont .
Oro gjorde mig sömnlös igår natt .
Torka dina tårar .
Djur kan inte särskilja mellan sant och falskt .
François , är denna din ?
Du skall observera trafikreglerna .
Syrien heter " Suriyah " på Arabiska .
Dayxa är min hustrus syster .
Dayxa är min svägerska .
Tom är den perfekta fadern .
Han kan inte utläsa vad det står på pappret .
Av någon anledning fungerade inte mikrofonen tidigare .
Var ser du tecknad film någonstans ?
Hon är en seriös person .
Jordskalvet skakade husen .
Jordbävningen skakade husen .
Jag håller på att dra ner på sötsaker .
Tuppen gal .
Han säger " kukeliku " .
Vad heter han nu igen ?
Han betedde sig som han borde .
Det var en obeskrivlig situation .
Hur som helst .
Var träffade ni varandra ?
Vi skulle i alla fall kunna försöka .
Mannen klagar , eftersom hunden skäller .
Eller är det tvärtom ?
Jag måste erkänna : jag ljög .
Om du vill prata så prata .
Behöver ni dricka vin ?
Mannen erkände slutligen vad han hade gjort .
Mannen erkände äntligen vad han hade gjort .
Mannen erkände till slut vad han hade gjort .
Delfinen är ett mycket intelligent djur .
Mannen erkände till sist vad han hade gjort .
Har posten kommit än ?
Han bor i den herrgården .
Han röstar alltid på Alliansen .
De är allierade .
Jag observerade att hans händer var ostadiga .
" Fina fisken " är ett exempel på svensk allitteration .
Ingen av oss vill gifta sig .
Hon är väldigt allmänbildad .
Våra föreläsningar är alltid öppna för allmänheten .
Vi måste komma på ett sätt att få den här maskinen att fungera under vatten .
Finns det några frågor av allmänintresse ?
Han är allmänläkare .
Det spelas inte mycket fotboll där .
De slog upp ett tält på en allmänning .
Jag vill gå med dig .
Jag älskar Lauries hår .
Vad gör du allra helst ?
Han tecknar en allriskförsäkring .
Där erbjöds allsköns aktiviteter .
Gud är allsmäktig .
De stämde upp i allsång .
På lördag är det allsångskväll .
Vem är allsångsledare i år ?
Allting har ett pris , det goda visar sig vara dyrare än det onda .
Vi tömmer förrådet allteftersom .
Tom stör Mary .
Det vet du inte .
Han har alltid varit vår alltiallo .
Han menar allvar .
Han såg väldigt allvarlig ut .
Det var en allvarsfylld tillställning .
Han tror sig vara allvetande .
Hon är en riktig allvetare .
Han köpte ett par allvädersstövlar .
Jag är en allätare .
En aln motsvarar femtionio komma trettioåtta centimeter .
Han föll ned i ett alnsbrett hål .
Han bor i en liten alpby i Österrike .
Alpfloran är mycket speciell .
Han tycker i en princip om alla alpina sporter .
Båten lade till nära kusten .
Vad vill du göra i framtiden ?
Han har alzheimer .
Vi pratade om diverse olika ämne .
Det hela utfördes på ett mycket amatörmässigt sätt .
Han är amatörskådespelare .
Ambassadbyggnaden är omgiven av höga stängsel .
Ambitionsnivån är hög .
Hon är den ambivalentaste människan jag känner .
Han fick åka ambulans till akuten .
Han fördes med ambulansflyg till Umeå .
Han arbetar som ambulanssjukvårdare .
Han utgör en del av ett ambulerande teatersällskap .
Hon är amfetaminmissbrukare .
Han är anhängare av amoralismen .
Hans amorbåge är helt perfekt .
Hur mycket amorterar ni på lånen ?
Snälla sänk volymen lite till .
Tom dödade Mary .
Tatoeba var tillfälligt otillgängligt .
Rädsla är skadligare än ett vasst svärd .
Kyoto är inte lika stort som Osaka .
Jag spelar volleyboll på stranden .
Jag är på stranden och spelar volleyboll .
Den här stanken får ju en att kväljas .
Jag förstår inte min klasskamrats kantonesiska .
Han tvingades amputera ena armen .
Han har amputerat bort ena benet .
Han har amputerat bort båda benen .
Hon slog an en ton på gitarren .
Han gick av och an i rummet .
Går han alltid an så där ?
Jag anade väl det .
Jag anade att någonting var på gång .
Han går på anabola .
Han är analfabet .
Har provet analyserats än ?
Vad är din analys ?
Vi bedömer också analysförmåga .
Han försöker anamma deras traditioner .
Han kan ingenting om anatomi .
En and simmade i vassen .
Några änder simmade i vassen .
Glöm inte att andas .
Hur stor andel får jag ?
Han förstod inte bokens andemening .
Hon blir andfådd av att gå upp för en trappa om tio trappsteg bara .
Han har andningsbesvär .
Lungan är ett andningsorgan .
Han gör aldrig andningspauser när han pratar .
Jag har vissa andningssvårigheter .
Han har långa andningsuppehåll nattetid .
Andra delen av boken var betydligt mycket bättre , tycker jag .
Hon bor i en andrahandslägenhet .
Förra månaden fick hon till slut ett förstahandskontrakt .
Vad heter du i andranamn ?
Har du något andranamn ?
Han hamnade på andraplats .
En andraplats är inte så dåligt heller .
Hennes andraspråk är franska .
Tar du andrastämman ?
Han är andratenor .
Alla andraårselever samlas utanför musiksalen .
Han är andretenor .
Han har ett väldigt androgynt utseende .
Morfar berättar gärna anekdoter .
Anfall är bästa försvar .
Du ska hålla ett anförande på minst fem minuter .
Jag vet inte vem jag kan anförtro detta åt .
Vem skulle anförtro honom någonting ?
Angav du källan till inkomsten ?
Det angav han inte .
Hans granne angav honom .
Han verkade väldigt angelägen när jag träffade honom sist .
Detta är en anglicism .
De angrep fienden i gryningen .
Personangrepp är inte tillåtna i forumet .
Vi tolererar inte personangrepp i kommentarsfälten .
Liisa är så försjunken i sin bok att hon inte ser eller hör någonting .
Norge och Sverige är angränsande länder .
Norge angränsar Sverige .
Det angår inte dig .
Vad angår det ?
Det går verkligen inte an .
Angående morgondagens möte : jag kommer inte att kunna infinna mig .
Nästa anhalt : Stockholm .
De anhöll en misstänkt i går .
Han anhöll om ett glas vatten .
Hans anhållan avslogs .
Kristendomen har många anhängare .
En anhörig identifierade kroppen .
Han har inga anhöriga .
Han är emot anhöriginvandring .
Han tittar gärna på animerad film .
Den där färgen var en aning bättre .
Hon har ingen aning om vad vi har planerat .
Han går som en anka .
Jag skulle önska mig att jag kunde uttrycka mig säkert , tydligt , vänligt och anpassat till situationen .
Liisa är så försjunken i sin bok att hon varken ser eller hör någonting annat .
Jag kan inte längre lita på dig .
Jag kan inte lita på dig längre .
Katten på bordet sover .
Misslyckandet fick Liisa att skämmas .
François , är detta ditt ?
Låt mig veta när du är klar !
Utan mig skulle du klara dig mycket bättre .
Körsbären blomstrar i april .
Det är klokt att spara för sämre tider .
Skruva ner tv : n .
Om jag ska säga sanningen minns jag ingenting jag sa i går .
Den kalla vinden plågade luffaren fruktansvärt .
Problemlösningen går framåt i snigelfart .
Min morbror bor i New York City .
Sjung ut !
Ut med språket !
De kom med vänner och fränder .
Jag blir inte klok på det .
Jag är utledsen på det .
Om det blir några svårigheter , ring mig !
Jag är urless på det .
Jag är utled på det .
Det här landet är en ankdamm .
Jag blir så trött på den här ankdammsdebatten .
Hon hade på sig en ankellång , röd klänning .
I går köpte jag tio nya par ankelsockor .
Vad anklagar du mig för ?
Det där är en väldigt allvarlig anklagelse .
Förslaget väckte stor anklang .
Förslaget vann stor anklang .
Han anknyter alltid till sin barndom i sina böcker .
Han äter alltid frukt som blivit ankommen .
När är deras beräknade ankomst ?
Vi möter er i ankomsthallen .
Ankomsttiden sköts upp tio minuter .
Han har mycket mjuka anletsdrag .
Vill du anlita mig ?
Vi måste anlita ett proffs .
Det är dyrt att anlita en advokat .
Tåget anlände en timme försenat .
Sista anmälningsdag är nästa fredag .
Har du skickat in din anmälan än ?
Anmälningsavgiften ligger på femtio kronor .
Du har anmälningsplikt .
Du är anmälningsskyldig .
Anmälningstiden har gått ut .
Måste du anmärka på allting ?
Huset var inte särskilt anmärkningsvärt .
Jag äter med händerna .
Informationen är hämtat ur de kinesiska annalerna .
Han är en mycket känd annalist .
Vi går någon annanstans och pratar .
Han satte in en annons i tidningen .
Med tidningen kom ett annonsblad .
Metro är en annonsfinansierad gratistidning .
Det råder annonsförbud här .
De har enorma annonsintäkter .
Din order har annullerats .
Han vill vara anonym .
Jag anar ugglor i mossen .
Detta hus har anor från 1800-talets slut .
Hon lider av anorexi .
Hon lider av anorexia .
Det är lika bra att anpassa sig .
Jag är anpassbar .
Hann du till bussen i morse ?
Hann du med tåget ?
Han går så fort att jag inte hänger med .
Hinner du komma på torsdag ?
Han hann .
Glöm inte att ta med dig en penna .
Stängde du av datorn när du gick hemifrån ?
Slår du på radion åt mig ?
Skruva upp volymen , är du snäll .
Vi hinner inte det i dag .
Vi får spara det tills i morgon .
Du är en bra bit på vägen .
Ingen har påstått det heller .
Är du på dåligt humör , eller ?
Nu ligger du illa till .
På vilken hylla ligger den ?
Fortsätt rakt fram och sväng sedan till höger .
Har du testat att starta om datorn ?
En omstart eller två brukar lösa de flesta datorproblem .
Bussen går om fem minuter .
Flyget avgår om fem minuter .
Tåget avgår om fem minuter .
Någon hade skräpat ned i trapphuset .
Kärlek och hosta kan inte döljas .
Jag fick lära mig den hårda vägen att det inte är klokt att köra bil när man är full .
Vad kostar denna penna ?
Jag har inte förstått .
Jag tror inte att de kommer att acceptera dessa villkor .
Min mage kurrar .
Jag är inte döv .
Vår plan har många fördelar .
Den här gamla fisken smakar konstigt
Jag har inte ätit något sedan i går .
De är lärare .
Hon är gift med en utlänning .
Ert rum är 504 : fem , noll , fyra .
Tom och Mary dricker ofta sitt morgonkaffe på verandan .
Du borde se den här filmen om du får chansen .
Jag minns detta ord .
Rum femhundrafyra är ert : femma , nolla , fyra .
Det har slutat att regna .
Finns det en bank nära stationen ?
Vad kostar den här kulspetspennan ?
Vad kostar denna kulspetspenna ?
Han krävde att hans lön skulle höjas .
Var på din vakt .
Höll ett öga öppet .
Jag minns det här ordet .
Eftersom jag inte hade varit länge i Tokyo , går jag ofta vilse .
Finns det någon bank nära stationen ?
Jag kommer ihåg det här ordet .
Det har slutat regna .
Han krävde en löneförhöjning .
Han krävde en lönehöjning .
Hon krävde en löneförhöjning .
Hon krävde en lönehöjning .
Kan du komma hit ett tag ?
Det kalla vädret fortsatte i tre veckor .
Han hade ett stort hus och två bilar .
Tom hade en benägenhet att titta bort när han blev tilltalad .
I alla språk finns det talesätt , fraser , idiom och ordspråk som inte kan översättas ordagrant .
De har inga barn , så vitt jag vet .
Den här föreningen grundades för etthundraelva år sedan .
I morse var jag uppe väldigt tidigt .
I morse var jag i farten väldigt tidigt .
Hur intressant !
Den här staden är tråkig .
Den här staden är död .
Troligen misslyckas han .
Han slängde många brev i papperskorgen .
Hon slängde många brev i papperskorgen .
Troligen misslyckas hon .
Du måste vara en idiot !
Priserna föll plötsligt .
I de flesta fall likställs modernisering med västernisering .
Han föregick med gott exempel .
" Vad är det här ? "
" Det är en persika . "
Egentligen ville vi gå på bio i lördags , men vi ångrade oss och stannade hemma .
Vad tänker du på just nu ?
Tvillingbröderna är lika som bär .
Vilken tid avgår bussen till flygplatsen ?
Vi firade hans födelsedag .
Hans hjälp kom i grevens tid .
Lådan är så lätt att den kan bäras av ett barn .
Sitter det en katt på bordet ?
När fadern kom hem , tittade jag på tv .
Hästen har fyra ben och snubblar ibland ändå .
Jag behöver ett frimärke .
Vi måste skjuta upp vår avresa .
Eftersom jag hade träffat honom en gång förut , kände jag igen honom direkt .
God afton , hur mår du ?
Jag står inte ut att bli störd i mitt arbete .
Ut ur mitt hus !
Han sökte i sin väska efter bilnyckeln .
Låt oss hoppas att hon kommer .
Jag spelar en timmes tennis varje dag .
Taket på mitt hus är rött .
Idag har jag hämtat min fyra år gamla brorson från dagis .
Hon är fem år gammal .
Jag vill sova lite längre .
Jag skulle vilja sova lite längre .
Han gifte sig med en skådespelerska .
Han gifte sig med en viss skådespelerska .
Han gifte sig med en viss skådespelare .
Hon gifte sig med en viss skådespelerska .
Hon gifte sig med en viss skådespelare .
Jag spelar tennis en timme om dagen .
Eftersom jag hade träffat honom en gång innan , kände jag genast igen honom .
Han är anpassningsbar .
Han är flexibel .
Människans anpassningsförmåga är unik .
Hon har vissa anpassningsproblem .
Han har köpt en anrik gård på landet .
Här anrikar man malm .
Vi har anropat förstärkning .
Han ansade skägget .
Grannen stod och ansade häcken .
Jag anser att det är onödigt .
Hon är en mycket ansedd konstnär .
Det skadade hans anseende .
Han köpte en ansenlig mängd råsocker .
Han har rena ansiktsdrag .
Alla i familjen har samma ansiktsform .
Han har gjort en ansiktslyftning .
Du skulle ha sett hans ansiktsuttryck .
Tycker du om ansjovis ?
Vilken anskrämlig soffa .
Har du anslutit HDMI-kabeln ?
Vi tar en anslutningsbuss till flygplatsen .
Vad anspelar du på ?
Du anstränger dig inte ens .
Detta är ett mycket ansträngande arbete .
Han såg ansträngd ut .
Hon hade ett ansträngt leende på läpparna .
Vi gör en sista ansträngning .
I höstas anställde vi fem nya medarbetare .
Är du anställd här ?
Har du fast anställning ?
I morgon ska jag på anställningsintervju .
Hur gick anställningsintervjun ?
Förslaget väckte anstöt .
Vem ansvarar för det här ?
Hon är ansvarsfull .
Han tar hand om ansvarsfördelningen .
Han ansökte om visum .
Har du ansökt om studiebidrag ?
Först måste du fylla i en ansökningsblankett .
Sista ansökningsdag är i övermorgon .
Nästa ansökningstillfälle är till hösten .
De antog förslaget .
Förslaget antogs .
Hans ansikte antog en lätt grön färg .
Det ska du inte anta .
Antagligen är det så .
Har antagningsbeskedet kommit än ?
Först måste du göra ett antagningsprov .
Han antastade henne .
Det är en oantastbar förmån .
Han är oantastbar .
Hon köpte ett nytt anteckningsblock .
Antecknar du ?
Han har skrivit en antibarbarus .
Han äter antibiotika .
Finns det något antikvariat här i närheten ?
Vilken färg har ditt hår ?
En tjej ringde mig .
Jag vet inte exakt när jag kommer att vara tillbaka .
Vad har du i din kasse ?
Jag pratar inte svenska .
Jag talar inte svenska .
Pratar du svenska ?
Jag pratar svenska .
Du kommer att tala svenska .
Ni ska tala svenska .
Ni kommer att tala svenska .
Ni kan förstå svenska .
Helga är ett svenskt namn .
Den som är född i Sverige är svensk .
" Är du svensk ? "
" Nej , schweizisk . "
" Är du svensk ? "
" Nej , jag är schweizisk . "
Hans fru är svenska .
Han tittade på en svensk film .
Jag tittade på en svensk film i går kväll .
Greta Garbo var en svensk skådespelare .
Antingen du eller jag måste göra det .
Har du installerat något antivirusprogram ?
Hans dikter publicerades i en antologi .
En antonym till synonym är antonym .
När är du anträffbar ?
Han var inte anträffbar .
Vad antyder du för något ?
Vad har papper för antändningstemperatur ?
Det här programmet är mycket användarvänligt .
Vilken användbar manick !
Vad har den för användningsområde ?
Aortan har spruckit .
Han spelar alltid apa .
Han apar efter alla andra hela tiden .
De utvisar apatiska barn .
I dag har jag tillryggalagt sex kilometer .
Vi använder apostlahästarna i stället .
Använd apostlahästarna !
När har apoteket öppet ?
Han har avlagt apotekarexamen .
Publiken applåderade .
Hunden apporterade .
Detta är bara ett approximativt värde .
Hon hade en aprikosfärgad klänning på sig .
Är detta ett aprilskämt ?
Vilket aprilväder det är i dag !
De träffades helt apropå .
Apropå lägenheter , vet du om dina föräldrar har hittat något nytt boende än ?
Jag har ingen aptit .
De spelade fyrhändigt .
De spelade à quatre mains .
De har köpt en ara .
Han kommer från en arbetarbakgrund .
Det råder arbetsbrist i landet .
Så här ser en typisk arbetsdag ut för mig .
Nu är ännu en arbetsdag över .
Vilken arbetsform föredrar ni ?
Vi måste komma överens om någon slags arbetsfördelning .
Du borde tala med din arbetsgivare .
Jag ska ut med en arbetskompis i morgon .
Arbetsledningen ignorerade förslaget .
Du har för lite arbetslivserfarenhet .
Han lever på arbetslöshetsersättning .
Vad säger arbetsmiljölagen ?
Han har hög arbetsmoral .
Du får se det som en arbetsmöjlighet .
Har filmen något arbetsnamn ?
Hur långt är ett vanligt arbetspass ?
Kan man få lite arbetsro här ?
Det är en gammal arbetsskada .
Hon har en gammal arbetsskada .
Det här arbetssättet passar mig inte .
I dag har jag varit i arbetstagen hela dagen .
Värst vad du är i arbetstagen .
En vanligt arbetsvecka börjar på måndag .
Argon är en ädelgas .
Är du arg på mig ?
Varför är du arg på mig ?
Var finns det en svensk ambassad ?
I går var det torsdag .
Jag vill ha en Toyota .
Vad har du för argument ?
Hon är duktig på att argumentera för sin sak .
Detta uttryck är arkaiskt .
Detta är en arkaism .
Han arkebuserades .
Han arbetar på ett arkitektkontor .
Hon deltog i en arkitekttävling .
Vi promenerade i staden och njöt av den vackra arkitekturen .
Han är mycket kunnig inom arkitekturhistoria .
Han har ingen riktig arkitektutbildning , men han jobbar ändå på landets finaste arkitektkontor .
Har du sökt i arkivet ?
Flera arkivalier har stulits .
Var snäll med din arma moder .
Armbandsur och armbandsklocka är två ord för en och samma sak .
Hon armbågade sig fram genom trängseln .
På Stockholms T-central måste man alltid armbåga sig fram .
Han skrapade upp armbågen .
Hon gjorde åttio armhävningar .
De gick i armkrok .
De gick arm i arm .
Du är under arrest .
Polisen har arresterat tre personer för lördagens inbrott .
Varför är du så arrogant ?
De har hittat tre nya arter i den här skogen .
Den här glassen innehåller massvis av artificiella ämnen .
Artikelförfattaren har bett om ursäkt för sin otillräckliga efterforskning i ämnet .
Just nu har tidningen en artikelserie om kvinnomisshandel .
Försök att artikulera mer när du sjunger .
Hon jobbar inom artistbranschen .
Han hoppas på en artistkarriär .
Han hoppas på en karriär som artist .
Hon använder sin hemort som sitt artistnamn .
Det ligger en artonhålsbana här i närheten .
Vittnen säger att vandalen var i artonårsåldern .
Hon arbetar på ett artotek .
Han har artros .
Jag kan inte stoppa blödningen .
Jag är 18 år gammal .
Jag talar inte tyska .
Jag är arton år gammal .
Språket är tungans musik .
Jag ska lära dig att spela schack .
Jag ska lära dig hur man spelar schack .
John är bra på schack .
John gillar schack .
Jag tycker om schack .
Ken slog mig på schack .
Vet du hur man spelar schack ?
Vad sägs om att spela schack i kväll ?
Jag vann över honom på schack .
Jag slog honom på schack .
Hur många olika pjäser är det i japanskt schack ?
Han har spelat schack sedan han gick på high school .
Har du några vapen ?
Vill du hänga ?
Vill ni hänga ?
Vill någon ha en öl ?
Ge mig inte den där blicken .
Tom försökte sälja sin gamla videobandspelare istället för att slänga den , men ingen köpte den , så det slutade med att han slängde den .
Tom sa att han inte var intresserad av Mary , men det verkade som att han alltid tittade åt den del av rummet som hon var i .
När jag läste till jurist sa mina lärare åt mig att aldrig ställa en fråga som jag inte visste svaret på .
När jag läste till advokat sa mina lärare åt mig att aldrig ställa en fråga som jag inte visste svaret på .
Din engelska är grammatiskt riktig , men ibland låter det du säger bara inte som något en modersmålstalare skulle säga .
Din engelska är grammatikalisk , men ibland låter det som du säger bara inte som någonting som en modersmålstalare skulle säga .
Han vande sig snart vid det kalla vädret .
Jag bodde i det här huset som barn .
Var är din skola ?
Dags att gå till skolan .
Var ligger din skola ?
Var ligger er skola ?
Det är dags att gå till skolan .
Krokodiler har vassa tänder .
En berusad man sov på bänken .
Jag bad Gud om en cykel , men jag insåg att det var inte hans metod .
Så jag stal en cykel och bad Gud om förlåtelse .
Busa inte !
Resultatet motsvarar inte mina förväntningar .
Hur klarar man av skolan när man knappt klarar av att ta sig dit ?
Jag kom ungefär klockan sex .
Ni behöver bara be om det .
Om du vill prata , prata då .
Om du vill prata , prata .
Jag vet bara vad Tom berättade för mig .
Jag ser honom ofta .
Att lära sig finska kräver tid .
Han råkade vara på samma tåg .
Vår tid är begränsad .
Han tömde sitt glas .
Han kom punktligt på utsatt tid .
Jag hörde det från en tillförlitlig källa .
Hur stavas det ?
Jag är inte det minsta orolig .
Ulster har minst förluster av alla boxare i ligan .
Jag är inte en pappersmugg .
Tom ser skräckslagen ut .
Ring brandkåren !
Jag kom vid sexsnåret .
Han har ett dåligt rykte bland sina studenter .
Vilket land kommer du ifrån ?
Hon säger att hon tycker om blommor .
Vi litar på honom .
Om det regnar i morgon , stannar vi hemma .
Jag kan inte hitta mitt bagage .
När de möter varandra , grälar de utan undantag .
Låt oss diskutera problemet med dem .
Var kan vi prata ostört ?
Var kan han hålla hus ?
Vad kan man göra åt det ?
Jag kan bara tala för mig själv .
Det bekymrar mig fortfarande .
Åt ni frukost ?
Jag är helt förvirrad .
Jag tvekar lite .
Känner ni dem ?
Känner du dem ?
Jag har anledning att anta att det inte är sant .
Det är svårt för människor att släppa gamla vanor .
Han kände medlidande med oss .
Det tog inte lång tid innan månen kom fram .
Tom kollade datumet .
Vad har du för bevis på att det var Tom som stal din mors halsband ?
Du har lättare för att komma ihåg saker än jag .
Jag vill att du går på mötet imorgon .
Du måste bli kvitt den där ovanan .
Du måste göra dig av med den där ovanan .
Hur kom du dit ?
Hur tog du dig dit ?
Hur ofta tvättar du dina jeans ?
Låt honom vänta ett ögonblick .
Låt honom vänta ett slag .
Glöm inte att det finns undantag .
Vilken blomma som helst går bra , så länge den är röd .
Tyvärr gick guiden fel .
Skrev du något i din dagbok idag ?
Tom ville inte tala med mig .
Tom ville inte prata med mig .
Häng din hatt på kroken .
Min katt hade ihjäl en ekorre .
Det här är ett mycket märkligt brev .
Det här är en mycket märklig bokstav .
Tom trodde att ingen var hemma .
Du behöver koppla av .
Är du lärare eller student ?
Den här maten är glutenfri .
Jag är allergisk mot gluten .
Var är rulltrappan upp ?
Mitt skosnöre fastnade i rulltrappan .
Det finns ingen regel utan undantag .
Jag håller inte med .
Han ser riktigt lycklig ut .
Vet du inte vem jag är ?
Vet ni inte vem jag är ?
Känner du inte igen Tom ?
Känner ni inte igen Tom ?
Ta reda på vad Tom vill .
Har du varit i Boston ?
Har ni varit i Boston ?
Har du hittat någonting ?
Har ni hittat någonting ?
Har du hört från Tom ?
Har ni hört från Tom ?
Han är flytande på Engelska .
Hur löste sig allt ?
Hur gick det med allt ?
Hur hamnade du här ?
Hur hamnade ni här ?
Hur kom du in hit ?
Hur kom ni in hit ?
Hur tog du dig in hit ?
Hur tog ni er in hit ?
Hur tror du att jag känner ?
Hur tror ni att jag känner ?
Hur tror du att jag känner mig ?
Hur tror ni att jag känner mig ?
Hur är ditt liv som gift ?
Hur är ert liv som gifta ?
Jag kan inte knäcka den här koden .
Jag kan inte ändra på vem jag är .
Jag kan inte göra det just nu .
Jag kan inte göra det längre .
Jag kan inte göra det här längre .
Jag kan inte låta dig göra det .
Jag kan inte låta er göra det .
Jag kan inte riktigt minnas .
Jag står inte ut med sjukhus .
Jag behövde inte din hjälp .
Jag behövde inte er hjälp .
Alla djur är lika , men vissa djur är mer lika än andra .
Jag skrev ingenting .
Jag skrev inte någonting .
Jag känner mig inte särskilt lycklig .
Jag måste inte vara här .
Jag tycker om inte den här platsen .
Jag gillar inte den här platsen .
Jag tycker inte om det här stället .
Jag gillar inte det här stället .
Jag fick ett F i kemi .
Jag har en till fråga .
Jag har en annan fråga .
De två försökte växelvis .
De två försökte ena efter den andra .
De köpte en ny dammsugare .
De har köpt en ny dammsugare .
De skulle köpa en ny dammsugare .
De ska köpa en ny dammsugare .
De kommer att köpa en ny dammsugare .
De kommer att ha köpt en ny dammsugare .
De skulle ha köpt en ny dammsugare .
De hade köpt en ny dammsugare .
De ska ha köpt en ny dammsugare .
Jag är homosexuell .
Kylskåpet är helt tomt .
Blir du inte trött i ögonen av att sitta framför en skärm hela dagarna ?
Har du kollat om vi har något bröd i frysen ?
Hittade du det du sökte efter ?
Han hittade inte det han sökte efter .
Han hittade inte det , som han sökte efter .
Är ugnen påsatt ?
Hur många grader ska ugnen stå på ?
Vilken temperatur ska ugnen stå på ?
Sitter du nu ?
Var bor du nu ?
Var bor ni nu ?
Var bor du just nu ?
Var bor ni just nu ?
Han fann inte det , som han sökte efter .
Han fann inte det han sökte efter .
Han respekterar inte mig .
Du måste respektera att han har en annan åsikt .
Jag uppskattar din ärlighet .
Det är ingenting som jag fäster någon vikt vid .
Han fäster stort avseende vid sådana saker .
Han har köpt ett bananfodral .
Det svider .
Det svider riktigt mycket .
Det svider till , men sedan går det över .
Det var ett svidande nederlag .
Hon staplade böckerna i en hög trave .
Hon backade in i en trave böcker .
Just nu har vi ett specialerbjudande för studenter .
Hur många armar har en bläckfisk ?
De ska åka på solsemester .
De ska åka på skidsemester .
De ska spendera semestern i fjällen .
De har stuga i fjällen .
Vilka fjäll brukar ni åka till ?
Hans största hobby är fjällvandring .
Han fiskar i en fjällbäck .
Vattnet i fjällbäckar är kristallklart .
De badade i det kristallklara fjällbäcksvattnet .
Han fyllde på sin vattenflaska i en fjällbäck .
Vem äger dessa renar ?
De har renar i ett hägn .
Gården är inhägnad av ett halvmeterhögt staket .
Jag tycker också om engelska .
Det fanns få barn i rummet .
Ge mig din tröja .
Om du inte vill dit , så åker vi inte dit .
Ingen vill dit .
Han agerade snabbt och släckte elden .
De tittade på teve .
Kan jag gå hem nu ?
Kan jag åka hem nu ?
Får jag gå hem nu ?
Får jag åka hem nu ?
De tittade på tv .
Han flög till Paris .
De är gymnasieelever .
Min far var ett träd .
Spanska är hans modersmål .
Mitt födelseår är 1982 .
Polisen fortsatte sin undersökning .
Har du någonsin varit i Rom ?
Han reflekterade över hur snabbt tiden går .
Jag föddes den tjugoandra november nittonhundrafyrtioåtta .
Var parkerade du bilen ?
Jag glömde boken hemma .
Denna punkt är värd att betona .
Det låter bekant .
Som pensionär är jag nu min egen chef - äntligen .
Denna punkt förtjänar särskild emfas .
Arbetet pågår .
Jämfört med henne är jag mycket opraktiskt .
Har ni någonsin besökt Rom ?
Den äldsta av oss kallas Mikko .
Spanska är hennes modersmål .
Det ligger inte alldeles här i närheten , men inte så långt borta heller .
Kan jag köpa enbart linserna ?
Var han fallskärmsjägare ?
Jag skulle vilja byta plats .
Tycker du om sommaren ?
Jag är korean .
Tom och Mary avskyr varandra .
Det liknar en anka .
Jag vill att du kommer tillbaka nästa vecka .
Vi vill inte skrämma bort barnen .
Vi hinner inte i tid till mötet .
Du pratar så fort att jag inte förstår ett ord av vad du säger .
Han stoppade näsduken i sin ficka .
Hans hus ligger precis över gatan .
Hans kropp hittades aldrig .
Datorreparationen tog hela dagen .
Hon är för ung för att skaffa körkort .
Bilden kostar tio pund .
Jag kan inte komma i dag , och inte heller i morgon .
Det där är en pagoda .
Inrättningen måste skyddas .
Du har druckit tre koppar kaffe .
Han är inget helgon .
Jag hade aldrig kunnat gissa att Tom och Mary skulle bli kära i varandra .
Det fanns mycket som vi helt enkelt inte hade tid att göra .
Jag gick upp tidigt för att hinna med tåget .
Smaklökar är väldigt användbara .
Brottslingen landsförvisades .
Jag kan inte tänka mig något annat .
Förutom borgmästaren var många andra förnäma gäster närvarande .
Det är svårt att utföra uppgiften .
Hur lång tid tog det honom att skriva den här romanen ?
Studerar du kemi ?
Pluggar du kemi ?
Tom är en hemmaman .
Hans svar var kort och koncist .
Alla säger att han ser ut precis som sin far .
Den här maskinen går på elektricitet .
Jag vinner .
De andra barnen skrattade .
Jag blev kär i dig .
Jag förälskade mig i dig .
Berätta om ditt dagliga liv .
Tom kunde inte hitta någon att prata med .
Jag önskar att jag hade varit med dig då .
Berätta om ditt vardagsliv .
Berätta om din vardag .
Hur lång tid tog det honom att skriva denna roman ?
Jag kan inte tänka mig någonting annat .
Jag steg upp tidigt för att hinna med tåget .
Jag klev upp tidigt för att hinna med tåget .
Ni har druckit tre koppar kaffe .
Han stoppade näsduken i fickan .
Tycker du om sommar ?
Hon tror att hon vet bäst .
Gud skapade jorden på sex dagar .
De gratulerade honom till hans bröllop .
Filosofi är inte ett så svårt ämne som du tror .
Försök en gång till .
Jag gillar kaffe mer än svart te .
Lyssnar du ?
Jag vill köpa .
Det är en timmes promenad till stationen .
Jag vill skicka detta paket till Kanada .
Jag vill skicka det här paketet till Kanada .
Det du fick lära dig är fel .
Det ni fick lära er är fel .
Det kräver bara lite beslutsamhet .
Det säger du alltid .
Jag behöver lite hjälp .
Var inte så nyfiken !
Han bär kläder i kinesisk stil .
Han bär kinesiska kläder .
Tycker ni att jag är ful ?
Frågorna hänger ihop .
Frågorna går in i varandra .
Jag måste göra det här själv .
Jag måste göra detta själv .
Jag tjänade precis tre lax .
Jag behöver bara hitta Tom .
Jag låste dörren på framsidan .
Jag behöver verkligen din hjälp .
Jag behöver verkligen er hjälp .
Jag sträckte ut armarna .
Jag sträckte ut benen .
Jag tror att jag är utarbetad .
Jag tror att jag är överansträngd .
Jag tror att det är bäst att du går .
Jag trodde att jag hörde musik .
Jag trodde att jag såg ett spöke .
Jag trodde att jag var i tid .
Jag trodde att det var ett skämt .
Jag trodde att Tom erkände .
Jag trodde att vi kunde prata .
Jag trodde att du hatade Tom .
Jag trodde att du gillade Tom .
Jag trodde att du tyckte om Tom .
Jag trodde att du åkte hem .
Jag trodde att du gick hem .
Jag trodde att du skulle gilla det .
Jag trodde att du skulle gilla den .
Jag trodde att du skulle tycka om det .
Jag trodde att du skulle tycka om den .
Jag trodde att ni skulle gilla den .
Jag trodde att ni skulle gilla det .
Jag trodde att ni skulle tycka om den .
Jag trodde att ni skulle tycka om det .
Jag trodde att ni åkte hem .
Jag trodde att ni gick hem .
Jag skulle hjälpa dig om jag kunde .
Jag skulle hjälpa er om jag kunde .
Jag skulle vilja tro dig .
Jag skulle vilja tro er .
Jag skulle vilja låna den här .
Jag skulle vilja låna detta .
Jag skulle vilja följa med Tom .
Jag skulle vilja träffa Tom nu .
Jag skulle vilja prata med Tom .
Jag skulle vilja tala med Tom .
Var inte så nyfikna !
Han är nykterist .
Dörren stängs automatiskt .
Det fungerar inte .
Den fungerar inte .
Var är kvinnan ?
Jag dödade Gud .
Jag vill inte gå till jobbet idag .
Det var fullmåne igår .
När serveras frukost ?
Jag dödade en gud .
Försök att sätta dig in i mitt ställe !
Du bad om det .
En man tog sig in på plan mitt under matchen .
Har du städat skrivbordet ?
Ta bara ett djupt andetag .
Skriv under på den sprickade linjen .
Ta Tom till stationen .
Det måste finnas ett mönster .
Tom åt en tidig middag .
Tom kan visa dig runt .
Tom kan inte lämnas ensam .
Tom dödade ingen .
Tom dödade inte någon .
Tom begick inte självmord .
Tom tog inte självmord .
Tom nämnde inte Mary .
Tom nämnde inte det .
Tom har inget hem .
Tom tog tag i Marys hand .
Tom har aldrig haft ett jobb .
Tom satte av mot dörren .
Har du fört över filmen till USB-minnet ?
Ligger filmen på USB-minnet ?
Hur stort är USB-minnet ?
Han hittade en gammal diskett .
Bilderna ligger på en cd-skiva någonstans .
Sitter cd : n i cd-läsaren ?
Jag är en morgonfrisk person .
Jag är en sjusovare .
Hur står det till ?
Jag är Döden .
Vi såg barnet stiga på bussen .
Om det bara vore så lätt .
Var är flygplatsen ?
De gick hand i hand .
Jag är här som turist .
Med den här jackan kommer du inte att frysa .
Jag hörde det på radion .
Var ligger flygplatsen ?
Var finns det en flygplats ?
Jag dricker inte ert vatten .
Hon köper bröd .
Jag väljer inte .
Jag älskar ingen .
Jag älskar inte någon .
Du behövde pengar .
Du hade behov av pengar .
I går var det dåligt väder här .
Han har en bror och två systrar .
Han är för gammal för er .
Hon är för gammal för er .
Tom är inte redo att ta emot gäster än .
Tom är inte redo att ta emot främmande än .
Tom var bara ett av Marys många fosterbarn .
Tom förberedde sig väl inför tentan .
Det var en skara människor i rummet .
Det var många människor i rummet .
Vems böcker är dessa ?
Vems böcker är de här ?
Vems böcker är det här ?
Vems böcker är detta ?
De är nöjda med det nya huset .
Jag är på väg till min systers bröllop .
Är det här din plats eller min ?
Är detta din eller min plats ?
Hos dig eller hos mig ?
Tom hade ingen anledning att bli arg .
Tom hade ingen anledning att vara arg .
Har du redan läst den här boken ?
Har du redan läst denna bok ?
Hunden är döende .
Tala långsammare .
Du förstår inte .
Ni förstår inte .
Denna produkt är tillverkad i Italien .
Den här produkten är tillverkad i Italien .
Ingen medicin kan bota denna sjukdom .
Ingen medicin kan bota den här sjukdomen .
Vi behöver dig .
Lyckan log mot henne .
Lyckan log mot honom .
Han hade mycket att göra .
Hon hade mycket att göra .
Du är vårt enda hopp .
Han gav mig ett exempel .
Kan du säga namnet på alla trädgårdens träd ?
Kan du säga namnet på alla träd i trädgården ?
Behöver du pengar ?
Jag åkte till flygplatsen för att träffa honom .
Jag åkte till flygplatsen för att möta upp honom .
De här tvillingarna är lika som bär .
Dessa tvillingar är lika som bär .
Mitt marsvin var min första flickvän .
Tom kommer att klara sig .
Tom döljer någonting .
Tom saknar ett finger .
Tom har timlön .
Tom är mycket fotogenisk .
Tom är blyg och feg .
Sverige är Skandinaviens största land .
Han dog i cancer .
Hon dog i cancer .
Utan honom är mitt liv tomt .
Utan henne är mitt liv tomt .
Detta är sant även i ditt fall .
Tom väntar på Mary .
Tom är inte rädd för dig .
Tom stirrade bara på Mary .
Tom sparkade omkull en stol .
Tom vet var Mary är .
Tom tittade på sin klocka .
Tom kollade på sin klocka .
Tom tittade på klockan .
Tom kollade på klockan .
Tom tittade på golvet .
Tom tittade i golvet .
Tom lyssnar aldrig på mig .
Tom såg honom aldrig igen .
Tom öppnade sin resväska .
Tom tog upp telefonen .
Jag har lite ont här .
Jag har ont här .
Hon köpte tre nya plektrum .
Hon köpte tre nya plektrer .
Spelar du med plektrum ?
Var la du plektrumet ?
Var la du plektret ?
Jag känner att jag sällan får någonting gjort .
Hur har din dag varit ?
Hade du några problem på vägen hit ?
Fungerar lokaltrafiken i dag ?
I går stod det helt still i lokaltrafiken .
Tog du bilen hit ?
Ta inte bilen , för parkeringen är stängd .
Lämna bilen hemma .
Tivolit är stängt under vinterhalvåret .
Den svenska vintern är mörk .
Popcorn är mitt favoritsnacks .
Popcorn är många gånger nyttigare än chips .
Hans största hobby är matlagning .
Försök att göra så liten åverkan som möjligt på väggar och golv .
Fick du mitt meddelande ?
Såg du inte att jag hade ringt ?
Han la ifrån sig mobilen när han var på stan .
Hur många watt är lampan på ?
Energilampor lönar sig i längden .
Var hittade du den här bilden ?
Läste du platsannonserna i tidningen i dag ?
Han platsar inte i laget .
Det vore verkligen på sin plats att hon bad om ursäkt .
Han har en platonisk kärlek till sin fru .
Hon har platinablont hår .
Han har plattfotsinlägg i sina skor .
Timme efter timme satt vi och lyssnade på hans plattheter .
En plattnäst kvinna kikade ut genom porten .
Hon samlar på plattänger .
Han köpte en reseplattång som fick plats i necessären .
De har parkerat uppe på platån .
Sverige duger inte för dem , så de firar alltid jul på playan .
Hon staplade sig fram i höga platåskor .
Det är en plausibel utkomst .
Det är en sannolik utkomst .
Fansen blev mycket besvikna när de märkte att stjärnan sjöng till playback .
Hon gör berlocker av plexiglas .
Han har pli på sin hund .
De har inte pli på sina barn .
Han är en pliktmänniska .
Han är en plikttrogen vän .
Plikttrogenhet är en egenskap som hon värdesätter högt .
Vem plingade i klockan ?
Hon plirade mot kameran .
Hon kisade mot kameran .
Jag öppnade dörren och såg ett par välbekanta , pliriga ögon .
En plirögd pojke vinkade till oss .
Han plitade ned några oläsbara bokstäver .
Han plitade ned en adress på ett solblekt papper .
Hon plitade ned sitt telefonnummer på baksidan av en gammal tidning .
De spelar plockepinn .
Han köpte plockgodis .
Han köpte lösviktsgodis .
Hon blir alltid dålig i magen av plockmat .
Äpplena är inte plockmogna än .
Har de plogat vägen än ?
Vi har en plogvall på garageuppfarten .
Plogbilen for nyss förbi på gatan .
Plogbilen åkte nyss förbi på gatan .
Han bär alltid plommonstop .
I trädgården står tre plommonträd .
Dagen till ära hade hon tagit på sig sin plommonfärgade aftonklänning .
Han dog av en brusten artär .
Om du inte lyssnar gör jag dig arvlös !
Hur stort är deras arvode ?
Du är inte arvsberättigad .
Hon har arytmibesvär .
Den där zombietjejen är uttryckligen döläcker .
Barnen tyckte att filmen var asbra .
Han var asberusad .
Hon lider av asbestos .
Tom är asexuell .
Hon låg tryckt mot den varma asfalten .
Asfalten var täckt med glassplitter från bilolyckan .
Välkommen till asfaltdjungeln !
Denna grusväg ska inom kort asfalteras .
De har asfalterat uppfarten .
Hon arbetar som asfaltläggare .
Du var asfull i går .
De asgarvade .
De asgarvar .
Alla asgarvar alltid åt hans skämt .
Hon är asiat .
Han la pengarna i en ask .
Jag är askblond .
Han är asket .
Han lever ett asketliv .
Hon är asocial .
Du var aspackad i går .
De finns många aspekter att ta hänsyn till .
Förra sommaren var himlen oföränderligt grå .
Det är många aspiranter på den här tjänsten .
Han aspirerar på chefspositionen .
Glöm inte att aspirera konsonanterna k , p och t när du talar svenska .
På finska aspirerar man inte konsonanterna k , p och t .
Han darrade som ett asplöv .
Kan jag få lite assistans här ?
Hon har assisterat oss i köket .
Den associationen får du stå för själv .
Det är din association och inte min .
Vad associerar du den här låten med ?
Han associerade den värma sommarvinden med frihet .
I en rimtävling gills inte assonanser .
Dessa är betygsatta på en hundragradig skala .
De vet inte hur en asterisk används .
Jag är astigmatiker .
Hon har astma .
Han fick ett astmaanfall .
Han fick en astmaattack .
Har du någon astmamedicin ?
Hon är astmatiker .
Han är astronaut .
Politikerna höll fester för astronomiska summor .
Det är inget konstigt att rymdprojekt kostar astronomiska summor pengar .
Spela på a-strängen .
Hennes konst präglas av en genomgående assymetri .
Hon målade assymetriska former på ett papper .
Gamar är asätare .
Han är ateist .
Detta är en ateistisk förening .
Han sitter i sin ateljé .
Klänningen är ateljésydd .
Han är atlet .
Ballongen svävade högt uppe i atmosfären .
Det var riktigt bra atmosfär på festen .
Attack är bästa försvar .
Östra flygeln är under attack .
Att-bisatser föregås ibland av kommatecken .
Jag gillar inte din attityd .
Hon har en förgräslig attityd .
Detta är helt och hållet en attitydfråga .
Vi behöver en attitydförändring i denna fråga .
De genomförde en attitydundersökning .
Ljus attraherar småkryp .
Småkryp attraheras av ljus .
Han är en mycket attraktiv man .
De fann diverse attrapper i mannens lägenhet .
Hon studerar audiologi .
Hon är audionom .
På denna skola utnyttjas många audiovisuella hjälpmedel i undervisningen .
Deras konsert planeras bli en audivisuell upplevelse .
Deras konsert planeras bli en audiovisuell upplevelse .
Hennes audition gick inte bra .
Han har bra auditivt minne .
Han har bra hörselminne .
Jag ska sälja mina gamla böcker på aktion .
Boken auktionerades ut för femhundraåttio kronor .
Hon arbetar som auktionsutropare .
Använd endast auktoritativa källor .
Han vill inte underställa sig auktoriteter .
Ö , ö , höö .
Det kan inte undvikas .
Haren springer i trädgården .
På grund av sjukdom kunde jag inte delta vid mötet .
På grund av sjukdom kunde jag inte delta på mötet .
Det går inte alltid som man vill .
Det går sällan som man vill .
Det är inte alltid lätt .
Hur svårt ska det vara ?
Det är bara att bita ihop .
Bit ihop nu !
Det är bara tre veckor kvar .
Kämpa på !
Hur ska man svara på den här frågan ?
Svaret på den här frågan finns inte i häftet .
Jag är fullständigt ointresserad av det här .
Utan intresse är det svårt att få motivation .
För motivation krävs ofta intresse .
Du har helt rätt .
Ni behöver bara be om den .
Nyheten om de två företagens sammanslagning kom ut igår .
Med några väl valda ord välkomnade han gästerna .
Hon invaldes i styrelsen .
Hon har selektiv hörsel .
Här finns det verkligen att välja och vraka bland .
Det här är min häst .
Detta är min häst .
Det är min häst .
Hästen är min .
Min pappa tog oss till djurparken igår .
På grund av sjukdom kunde jag inte delta i mötet .
Han föll huvudstupa i vattnet .
Hennes dotter har alla förutsättningar för att bli en bra lärare .
Åt du frukost ?
Det är dags att öppna den tredje garderoben .
Detta kan vara korrekt .
En av dem slog mig i ryggen .
Vad fan gör du här ?
Jag har tillräckligt med pengar för att köpa en bil .
Ditt rum är dubbelt så stort som mitt .
Jag ringde inte honom eftersom jag hade en förkylning .
Vi tar kreditkort .
De förklarade sig oskyldiga .
Ett bi surrar .
Det största sovrummet har söderläge .
Det största sovrummet vetter mot söder .
Har du varit på Koreahalvön ?
Jag såg bilen köra på en man .
Den här boken behandlar Kina .
Mitt rum vetter mot öst .
Faktum är att han inte håller med mig .
Faktum är att han är troende .
Soldaterna är döda .
Torka byxorna på elementet .
Tom har aldrig ätit rått hästkött .
Olyckligtvis släppte Tom ut katten ur säcken .
Vi såg något vitt i mörkret .
Tom tycker inte om den här färgen .
Tom kunde knappt gå .
Jag gick längs huvudgatan .
Jag kan inte fatta att vi äntligen klarade det .
Det är inte tillåtet för kvinnor att köra bil i Saudiarabien .
Det finns blott ett alternativ .
Han är säker på att det är curry .
Hur bred är den här vägen ?
Jag uppfattade inte riktigt namnet på den där designern .
Flyger du ofta ?
Flyger ni ofta ?
Får den här lådan plats i skåpbilen ?
Den här hunden är min .
Sådant kan hända då och då .
Hon kunde inte hindra sin dotter från att gå ut .
Jag köpte många böcker .
Jag köpte en massa böcker .
Förlåååt .
Jag kunde inte sova i går kväll , så jag försov mig .
Hihi !
Han är längre än sin bror .
Han är längre än sin lillebror .
Han vet bättre än att gifta sig med henne .
Jag älskar Kalifornien .
Jag arbetade på en bondgård .
Musikern är känd i utlandet såväl som i Japan .
Hon lever på grönsaker och råris .
Jag kokar fortfarande råriset .
Jag har ätit svartrissoppa tre gånger på en dag !
Luften är fuktig .
Chongqing är en kuperad stad med slingrande vägar .
Ingen vet säkert hur många människor som dog .
Hon har inga barn .
Hon har små bröst , men jag har inget emot det .
Jag känner mig lättare än luft .
Vill du gå någon annanstans ?
Hans tal fångade vår uppmärksamhet .
Jag glömde ditt paraply på bussen .
Han låter den här pistolen vara laddad .
Min far , farfar , farfars far och farfars farfar hade alla samma namn som jag .
Toms farfar och Marys farfar slogs tillsammans i andra världskriget .
Toms farfar och Marys morfar slogs tillsammans i andra världskriget .
Toms morfar och Marys farfar slogs tillsammans i andra världskriget .
Toms morfar och Marys morfar slogs tillsammans i andra världskriget .
Vi döpte min son efter min farfar .
Vi döpte min son efter min morfar .
Spädbarnet döptes till Alfred efter sin farfar .
Spädbarnet döptes till Alfred efter sin morfar .
Tom tvivlar inte på Marys förmåga att utföra jobbet .
Bill , ring mig ikväll .
Känner du till kabuki ?
Första steget är det jobbigaste .
Jag tycker inte om honom , för han är slug som en räv .
Han är en slug räv .
Han har kommit att se ut att vara en rävaktig premiärminister som utnyttjar makten i sitt ämbete till fullo för egen vinning .
Tunnelbanan går under jord .
Det är billigt att åka tunnelbana i Peking .
Jag tvivlar på att Tom är glad .
Jag tvivlar på att Tom är lycklig .
Sitter du här och ugglar nu igen ?
Vi måste undersöka denna fråga i förväg .
Jag är så upptagen att jag inte kan hjälpa dig .
Jag skulle aldrig säga något sådant .
Tycker du att jag är ful ?
De älskar varandra väldigt mycket .
Jag läste ut boken i går kväll .
Det går inte att förutsäga vad som kommer hända nästa år .
Jag är inte galen .
Jag gillar inte huset .
Bröd bakas i ugn .
Bröd bakas i en ugn .
Det var en av mitt livs mest makalösa upplevelser .
Den tycker om att röka tobak .
Det tycker om att röka tobak .
Jag åkte till Italien för andra gången 1980 .
Kontrasten mellan himlen och berget är slående .
Tom dyker oftast upp i tid .
När såg du senast Tom ?
Kom ner så snart som möjligt .
Tom har aldrig sett Mary så arg .
Stormen sänkte temperaturen .
Jag har inte druckit kaffe än .
De övertalade mig att stanna ett tag till .
Jag är rädd för vilda djur .
Jag ska ta den jäveln .
Mary har all anledning att vara nöjd .
Varför frågar du mig ?
Vi spelar schack .
Jag har redan tagit fyra av hans pjäser .
Gruppen springer på stranden .
Gör dig av med pistolen .
Jobbar du fortfarande med Tom ?
Arbetar du fortfarande med Tom ?
Jag väntar på att affärens ska öppna .
Fastän de ser ut som det är Carlos och Juan inte enäggstvillingar , bara bröder .
Jag bestämde mig för att jag inte ville ha mer med Tom att göra .
Hon är lång och smal .
Han lovade mig att vara mer försiktig i framtiden .
Hantverkaren lovade att komma nästa dag .
Plutonium-239 har en halveringstid på 24 100 år .
Tom undrade varför Mary var så sen .
Jag är egyptier .
Jag var nära att dö av en hjärtattack .
Jag hittade en fin lägenhet åt honom .
Tom vill att Mary ska träffa hans mor .
Finns du ?
Finns de ?
Var det här någon annans idé ?
Oavsett vad som händer kommer jag aldrig att ändra mig .
Det här vinet smakar gott .
Det här vinet är gott .
Varför skulle någon vilja göra det ?
Jag hörde någon skrika .
Jag stod en stund och tittade på avgasröret .
Kort hår passar henne verkligen .
Jag tänker skriva om våra parker och berg .
Kineserna vet inte att jag inte är mänsklig .
Vi stötte på dem vid bussterminalen .
Jag vill ha ett par handskar .
Hörde du klickljudet ?
Jag tror inte mina ögon .
Jag trodde inte mina ögon .
Jag trodde knappt mina ögon .
Han trodde inte sina ögon .
Det är alltid värt ett försök .
Jag minns hans ansikte , men jag kommer inte ihåg hans namn .
Han kommer alltid till klassträffarna .
Du måste passa din hund .
Jag tror du har rätt .
Jag tror att du har rätt .
Jag vet att du inte ville att Tom skulle åka in i fängelse .
Hennes namn är känt världen över .
Hans namn är känt världen över .
Jag är van vid att arbeta hårt .
Hörde du mig inte ?
I morgon är det samling i aulan .
Hon arbetar som au pair i Tyskland .
Han är australier .
Han är australiensisk .
Hon är australiensiska .
Han är australisk .
Detta är en autentisk källa .
Han är min favoritauteur .
Deras son har autism .
Deras son är autistisk .
Fotograferar du med autofokus ?
Kan jag få din autograf ?
Skulle jag kunna får din autograf ?
Det sker automatiskt .
Tillverkningen har automatiserats .
Han misstog bilens farthållare för autopilot .
Har du avaktiverat tjänsten ?
De avancerade nivåerna är riktigt svåra .
Jag vill avanmäla mig .
Har ni avbeställningsskydd ?
Vi har den perfekta avbetalningsplanen för dig .
Hon köpte den på avbetalning .
Hennes breda bak hade avbildats i form av ett rumpavtryck i soffan .
Knip av tråden med en avbitare .
De var tvungna att avblåsa matchen .
De var tvungna att blåsa av matchen .
Har du avbokat vårt bord ?
Varför avbryter du mig hela tiden ?
Kan jag få tala till punkt , utan att du avbryter mig ?
Vi ursäktar avbrottet .
Vi måste tyvärr avböja ert anbud .
De fick poängavdrag .
Resan måste avbeställas senast tjugofyra timmar innan avresa .
Det verkar som att den självrättfärdige tölpen äntligen är borta .
Hon stirrade in i hans tättsittande ögon .
Det här är ingen tävling .
Jag vandrar i ett töcken .
Jag har endast töckniga tankar inför framtiden .
Han är en tävlingsmänniska .
Det har börjat töa .
I dag är ännu en töig dag .
Ditt stora huvud töjer ut den .
Tröjan är ganska töjbar .
Tummis på det !
Det bidde bara en tumme av det hela .
Han har tummen mitt i handen .
Jag håller tummarna för dig .
Kan vi träffas på tumanhand ?
Han har en riktig tjurnacke .
Vad är han där för en tjomme ?
Tjosan hejsan !
Jag åkte aldrig fast .
Det visade sig att han visste allt om mig .
Tom och Mary har en mack ihop .
Jag köpte mackan på macken .
Tomten är inte till salu .
Russin är skrumpnade vindruvor .
Russin är torkade vindruvor .
Tom åt en handfull russin .
Du skulle ha sett henne .
Det är hälsosamt att vara galen .
Du gör mig förbannad !
Sex var inbjudna , pojken inkluderad .
Vad ska du göra ikväll ?
Det här trädet är inte ens i närheten av att vara det högsta i socknen .
Kan de se oss ?
Du har förlorat koncentrationsförmågan .
Tror du på spöken ?
Hon är mer vis än smart .
Han verkar inte ha vetat det .
Vad äter vi ikväll ?
Vad tänker du på ?
Den internationella konferensen skulle gå av stapeln i februari i år .
Festivalen kommer att gå av stapeln nästa vecka .
När bröt andra världskriget ut ?
Jag åker dit varje år .
Jag har aldrig varit hemma hos min farbror .
Jag har aldrig varit hemma hos min morbror .
Det är oartigt att peka på folk .
Jag kommer inte ihåg vilka artiklar jag har översatt och inte .
Han sprang för att komma i tid .
Jag köpte smörgåsen på macken .
Hon drog mig åt sidan .
Huset föll samman i ett jordskalv .
Huset föll samman i en jordbävning .
Ta min .
Ta mitt .
Tag min .
Tag mitt .
Låt mig gå !
Det är fullständigt omöjligt att ni åker till New York den här helgen .
Vi ses i morgon !
Skulle du kunna berätta hur man tar sig till stationen ?
Han fuskade på biologiprovet .
Han fuskade på biologitentan .
Han fuskade på biologitentamen .
Han sa att han inte vet .
Han sa att han inte visste .
Koste vad det kosta vill .
Hon är alltid väldigt artig .
Han bygger en bro .
Han sitter i isoleringscell .
Ingen får gå dit .
Han höll på att bli en känd sångare .
Vill du ha lite mer nötkött ?
Vad är lufttemperaturen idag ?
Säg någonting även om du inte vet rätt svar .
Han går upp tidigt .
Han stiger upp tidigt .
Jag tittade på henne .
Jag hoppas att få se renar under min resa till Sverige .
Tom borde ha varit här vid det här laget .
Tom sa att han ville komma bort från stan ett tag .
Tom sade att han ville komma bort från staden ett tag .
Var student har sin egen dator .
Varje student har sin egen dator .
Var elev har sin egen dator .
Varje elev har sin egen dator .
En förbipasserande filmade polisens våld med sin mobiltelefon .
Har du pojk- eller flickvän ?
Var träffade du hen ?
Har du pojk- eller flickvän ?
Var träffade du honom eller henne ?
Jag vill bara kunna besöka mina barn när jag så önskar .
Jag vill bara kunna besöka mina barn när jag vill .
Jag stannade hemma i går kväll för att kunna ta emot ditt samtal .
Har du någon hostmedicin ?
Har ni någon hostmedicin ?
Jag bryr mig inte om vad de säger .
Det rör mig inte i ryggen vad de säger .
Det rör mig inte i ryggen .
Flickan stirrade på dockan .
De blev mördade .
De mördades .
De var perfekta .
De var mina .
De var hjältar .
De var falska .
De vill ha mig .
De ville ha bevis .
De blev tokiga .
De litar på dig .
De började dansa .
De började skjuta .
De tog i hand .
De skakade hand .
De ser bra ut .
De ser förvirrade ut .
De gick ut .
Om du är upptagen nu kan jag ringa tillbaka till dig senare .
Tar ni det här kortet ?
Skyskrapan förväntas sjunka ner i myren .
Varför tror du att jag tänker på dig ?
Råttor förökar sig snabbt .
Var har hon köpt de här böckerna ?
Marknaden öppnar klockan nio på morgonen .
Jag trodde du var van vid att bo i husvagn .
Toms föräldrar bor i en gammal husvagn .
Han kopplade på husvagnen på sin bil .
Lite skit rensar magen .
" Kebabmorden " verkar ha lösts .
Årets icke-ord 2011 är " Kebabmord " .
Det är bara en teori .
Hur tung är er väska ?
Var snäll och glöm inte att skriva med stora bokstäver .
Var snäll och glöm inte att skriva med versaler .
Jag letar efter en man som ska bo här .
Jag tror inte att tv någonsin kommer att ersätta böcker .
Jag vill inte störa Tom .
Kan jag få tala med henne ?
Han beskrev olyckan i detalj .
Tro inte på henne , hon ljuger alltid .
Vi får inte många besökare här nere .
Om du tänker döda mig så vill jag veta varför .
Tom borde inte ha ätit så mycket .
Hur dags går nästa tåg till Tokyo ?
Min bror måste skriva en tentamen .
Jag tycker om att översätta dina meningar .
Jag är bög .
Min skrivare skriver bara ut i svartvitt .
Laserskrivare är generellt sett billigare i underhåll än bläckstråleskrivare
Fladdermusen är inte en fågel , utan ett däggdjur .
Han måste städa sitt rum .
Han borde ha vetat bättre .
Han kliver upp tidigt .
Hon tycker mycket om att gå på bio .
Vi måste vänta på honom .
Han sover som en bebis .
Njut av ögonblicket !
Jag känner mig lite svag idag .
Det var ett riktigt stort rum .
Hans ord sårade Meg .
Hon besökte sin man i fängelset .
Stäng dörren !
Det drar .
Jag tillbringade min semester utomlands .
Jag pantsatte min gitarr för att betala hyran .
Jag pantsatte min gitarr så att jag kunde betala hyran .
Polisen undersökte de misstänktas antecedentia .
Jag har inte kunnat gå till skolan på en vecka .
Jag har en dator .
Vänta här tills jag kommer tillbaka .
Jag värmer inte upp deras hus åt dem .
Tom kan inte göra någonting utan Marys hjälp .
Eleverna har tillgång till dessa datorer .
Hon har stora bröst .
Hungrig ?
Hon tillhör tennisklubben .
I detta land ser man överhuvudtaget ingen skillnad på arbetstid och fritid .
Skulle du kunna förklara hur man tar sig dit ?
När du är i Rom , bete dig som romarna .
Här är jag född och uppvuxen .
Fetma är en nationell epidemi .
Jag fick en massa myggbett .
Mamma var allt som oftast väldigt upptagen .
Varför är du så trött ?
Han är van vid att gå långa sträckor .
Jag vill inte leva .
Den här boken tillhör mig .
Tack för att du tröstade mig när jag var ledsen .
Denna teori kan jag inte acceptera .
Hon är på riktigt gott humör .
Jag kan inte tänka mig ett liv utan dig .
Jag flyttade till en ny lägenhet .
Arbeta inte för mycket .
Försöket misslyckades .
Tom försvann utan att lämna ett spår .
Klä på dig fort .
Klä på er fort .
Det är fyrtioåtta sjömän på skeppet .
Han drack direkt ur flaskan .
Hennes syster bor i Skottland .
Tom försvann utan ett spår .
Ju galnare , desto bättre .
Du måste ha tålamod .
Ni måste ha tålamod .
Tycker du om klassisk musik ?
Detta kan leda till otrevliga konsekvenser .
Det var dags att gå .
Kineserna är hårt arbetande människor .
Hur använder man ätpinnar ?
Vi har sett henne .
Hon har sönder något varje gång hon städar rummet .
Snabba er , ungar , annars missar ni skolbussen .
1891 blev Liliuokalani Hawaiis drottning .
Jag kunde inte somna .
Allt gick bra .
Det finns nästan inget syre i rummet .
Det här är mina byxor .
Det här företaget använder billig arbetskraft för att öka sina vinstmarginaler .
De bor i en liten by i England .
Två läsk till barnen och en kaffe , tack .
Hur många dagar gammal var jag när den här bilden togs ?
" Den gamle och havet " är en roman av Hemingway .
Det bodde en gubbe i det gamla huset .
Det bodde en gammal man i det gamla huset .
Det bodde en gammal gubbe i det gamla huset .
Gubben är blind på ena ögat .
Den gamle mannen är blind på ena ögat .
Du får prata hur mycket du vill .
Han lider av en svår sjukdom .
Tom är vänsterhänt , men han skriver med höger hand .
Jag skrev till honom av en helt annan anledning .
Tom kommer inte att döda någon annan .
Jag skulle vilja ha något att dricka .
Den här kameran är tillverkad i Tyskland .
Jag kompenserar för det nästa gång .
Han har hår på bröstet .
Hon är inte vackrare än deras mor .
Han rånade en gammal dam .
Max förklarade för Julia varför han inte kunde komma på hennes avskedsfest .
Det här är en väldigt tidsödande uppgift .
Jag vill verkligen inte lämna barnen ensamma nu .
Jo-Jo var en man som trodde att han var en ensamvarg .
Jag har alltid varit en ensamvarg .
Jag är något av en ensamvarg .
Tom vill inte prata med dig .
Hans rum är alltid i ordning .
Vi har åtminstone tak över huvudet .
Denna bok , som jag har läst två gånger , var en present från Peter .
Han var tyst av rädsla .
Tom dricker inte .
Hur många dagar var jag när den här bilden togs ?
Gillar du klassisk musik ?
Vad heter denna gata ?
Jag försöker bara tjäna en slant .
Fastän det låter märkligt är det sant det hon sade .
Hon hittade jobb som maskinskriverska .
Han känner inte mig .
Ibland förstår jag mig inte på honom .
Ibland förstår jag inte honom .
Ibland förstår jag honom inte .
De gjorde honom till klubbens ordförande .
Jag har bara sett det en gång .
Jag har bara sett den en gång .
Vad är klockan ?
Vad sägs om en kopp te ?
Vet du hur hans far dog ?
Han skadades allvarligt i trafikolyckan .
Var snäll och tänd lampan .
Men jag kan inte grilla grillspett !
Jag kan inte använda vänster hand på grund av gipset .
Den är tom.
Det är tomt .
Vilken lättnad !
Vilken relief !
Ge mig något att skriva på .
Ge mig något att signera .
De fångade rävar med fällor .
Något kommer att hända .
Jag känner det på mig .
Var någon annan frånvarande ?
Ungarna spelar Duck Hunt .
Barnen spelar Duck Hunt .
Jag var tvungen att överge min plan .
Jag vill att du kommer tillbaka till Boston .
Det är en encellig organism .
Detta var en skön känsla .
Hon ser vacker och frisk ut .
Din katt är tjock .
Er katt är tjock .
Hur snart måste jag vara tillbaka ?
Maten var hemsk , men jag har inte klagat .
Jag för dem till Kate .
Det är en skugga .
Hon är van vid att sitta .
Jag hoppas att det ska vara bra imorgon .
Företaget vill anställa 20 personer .
Tom kom hit för att be oss om hjälp .
Tom kom hit för att be om vår hjälp .
Tror och tror , det handlar snarare om övertygelse .
Vill du ha lift ?
Vill du ha skjuts ?
Det tog mig en halvtimme att lösa det här problemet .
Hon är nästan sextio år gammal .
Jag tänker så det knakar , men jag kan inte komma på hennes namn .
Våldet varade i två veckor .
Du är annorlunda .
Damer och herrar , välkomna ombord .
Tom känner inte att han kan lita på Mary .
Tom masserar sina knän .
Tom masserar hans knän .
Tom klagar nästan aldrig på någonting .
Hennes argument byggde inte på fakta .
Vill du gifta dig först eller skaffa barn först ?
Kan du höja volymen på radion litet ?
Jag trodde att valar är fiskar .
Tom dricker inte öl .
Jag såg månen ovanför taket .
Jag vill ha fem köttbullar .
Kan du skriva ner det ?
Kan jag ta ett meddelande ?
Han är inte min pappa .
Kan du skriva ned det ?
Vill du gifta dig eller skaffa barn först ?
Företaget vill anställa tjugo personer .
Jag hoppas att det är bra i morgon .
Det här var en skön känsla .
Någonting kommer att hända .
Jag känner det på mig .
Tom undrade om det Mary sa var sant .
Fastän det låter märkligt är det hon sade sant .
Tom häller upp ett glas mjölk .
Det blir tre euro .
Tom var gift på den tiden .
Jag var så lycklig på den tiden .
Tom kunde inte bestämma sig .
Vi trodde att hans hot bara var ett skämt .
Han får göra vad han vill med pengarna .
Han kan göra vad han vill med pengarna .
Jag träffade ingen på vägen hem .
Den här pojken är lat .
Tom behöver sannerligen inte mer pengar .
Det är inget skämt .
Hans otrevliga kommentarer spädde på dispyten .
Vilken underbar trädgård !
Målet var offside .
Jag har bott här hela mitt liv .
Tom låtsades inte höra Mary ropa hans namn .
Berätta för Tom vad du vill göra .
Jag är mördaren .
Jag kan simma bra .
Den här romanen är översatt från engelska .
Tom tänkte inte på det .
Det här är ett postkontor och det där är en bank .
När kan vi träffas igen ?
När kan vi ses igen ?
Hon är ungefär i min ålder .
Jag köpte den här kameran för 35 000 yen .
Vi har inget annat val .
En färsk undersökning visar att antalet rökare minskar .
Vad gjorde du med den här boken ?
Vad gjorde du av den där boken ?
Titta på pojken bredvid bilen .
Den här boken innehåller fyrtio fotografier .
Jag har ett tajt schema den här helgen .
Det var svalt och skönt , men nu börjar det bli kallt .
Frihetsgudinnan är symbolen för USA .
Jag kan inte engelska .
Jag önskar att jag vore ung igen .
Min mor sade åt mig att uppföra mig .
Han tycker om att spela tennis .
Jag vill lära mig att spela go .
Lär av kamrat Lei Feng .
Hon var på dåligt humör .
Jag vill inte sjunga , för jag är tondöv .
Han inser inte att han är tondöv .
Vem kan utföra det här arbetet ?
Elefanter är majestätiska djur .
Vem spelar huvudrollen ?
Väntar du på oss vid stationen ?
Väntar du på oss på stationen ?
Väntar ni på oss på stationen ?
Väntar ni på oss vid stationen ?
Kommer du att vänta på oss på stationen ?
Kommer du att vänta på oss vid stationen ?
Kommer ni att vänta på oss vid stationen ?
Kommer ni att vänta på oss på stationen ?
Han tog fram några mynt .
Han tog ut några mynt .
Det var just likt honom att komma för sent .
Jag ämnade att lyckas , men kunde inte .
Jag tvättade medan spädbarnet sov .
Kärnvapen är ett hot mot hela mänskligheten .
Hon gråter alltid när han är full .
Han gråter alltid när han är full .
Vi spelar ofta schack .
Du vet den där känslan ?
Svarta katter betyder otur .
Vad fattas dig ?
Du ser blek ut .
Du ser blek ut idag .
Vem upptäckte Amerika ?
Varför skär du upp frukterna ?
Ibland är det viktigt att fatta ett beslut snabbt .
Hon hade på sig en svart hatt .
Gråter du ofta ?
Du litar fullständigt på honom .
Ni litar fullständigt på honom .
Du dödade Tom .
Ni dödade Tom .
Asken , som jag hade hittat , var tom.
Jag tror att det är omöjligt att förneka detta faktum .
Tom överraskade Maria med en kyss .
Bröllopet sköts upp .
Nu eller aldrig .
Det skulle vara trevligt om jag kunde resa till Japan .
Han har två döttrar .
Du gjorde det mycket bra .
Det fattades bara !
Jag är ledsen att du fick vänta .
Han spelade piano .
Hon var klädd i svart .
Han förlorar aldrig hoppet .
Framför mitt hus finns en sjö .
Du är lat !
Ni är lata !
Vad tittar du på mig för ?
Vad tittar ni på mig för ?
Vill du att jag ska hålla ett öga på Tom åt dig ?
Hon var inte snabb nog .
Hon var inte tillräckligt snabb .
Det är tydligt att han är hemma .
Jag har matteläxa idag .
Är du redo att beställa nu ?
Är ni redo att beställa nu ?
Det här spelet är baserat på en roman .
Han studerade hur fåglar flyger .
Hitta katten .
Jag spelade fotboll igår .
Kvinnan är rik , men mannen är fattig .
Man kan inte stoppa tillbaka tandkräm i tuben .
Populisterna har vunnit .
Jag fick veta att det var svårt för henne att lösa det problemet .
Tåget bör vara i Osaka vid tio .
Den här medicinen kommer att bota din förkylning .
Vilket som .
Det är oviktigt .
Jag åkte flygplan till Kyushu .
Jag tycker inte om det .
Jag tycker inte om det där .
Jag gillar det inte .
Det besegrade laget lämnade så sakta planen .
Stick !
Vår bil är tre år äldre än er .
Vår bil är tre år äldre än din .
Vår bil är tre år äldre än era .
Vår bil är tre år äldre än dina .
Varför denna kalabalik ?
Han håller på att bli skallig .
Jag åkte till Kyushu med flygplan .
Det gjorde du mycket bra .
Föräldrarna försökte att avdramatisera barnets tandläkarbesök .
De promenerade längs avenyn .
De återvinner alla sina hushållsavfall .
De återvinner allt sitt hushållsavfall .
Han var mager och avfallen .
Det ligger en avfallsanläggning på andra sidan berget .
Han bodde i en avfallshög .
Vilken avfart ska jag ta ?
De svängde av på fel avfart .
Ni måste ha tagit fel avfart .
Är det nästa avfart vi ska ta ?
Har du avfettat alla maskindelar ?
Har vi något avfettningsmedel ?
De måste avfukta källaren .
Hon avfyrade ett skott i luften .
I morgon är det avfärd .
De avförde ärendet från dagordningen .
Han började hosta av alla avgaser .
Rummet fylldes av avgaser .
Bilen täcktes i ett avgasmoln .
Den här bilen har två avgasrör .
Nu tillkommer det nog inte fler avgifter .
Res inte med dem .
De har alltid så många dolda avgifter .
Han är inne på avgiftning .
Snart kommer också läsplattor att avgiftbeläggas .
Hon föll ned i en avgrund .
Det här stupet är avgrundsdjupt .
Hon gav ifrån sig ett avgrundsvrål .
Du måste avgränsa ditt forskningsområde ytterligare .
Flyget avgår om fyrtiofem minuter .
Han avgick efter sexskandalen .
Hon stoltserade med sitt avgångsbetyg .
Dagens match är avgörande .
Det blev ett snabbt avgörande .
Hon har skrivit en avhandling på traditionell kinesisk medicin .
Det har skett många avhopp på sistone .
De försöker att avhumanisera asylsökande , och vinner därigenom opinion .
Förra året avhystes en hyresgäst i huset här bredvid .
Hon medverkat i några mycket avhållna filmer .
Han är avhållsam .
De förespråkar avhållsamhet i alla sina former .
De hängde av sig ytterkläderna i hallen .
Vill du ha din avi per sms ?
Han är bara avis .
Han är bara avundsjuk .
De avisade bron med salt .
Jag kommer inte att behöva dig .
Jag kommer inte att behöva er .
Äta bör man , annars dör man .
Äta bör man , annars dör man .
Äta gör man , ändå dör man .
Undra vems bil det här är .
De steg ombord på flygplanet .
I början förstod jag inte varför .
Där fanns inte en kotte så långt ögat kunde nå .
Där fanns inte en levande själ så långt ögat kunde nå .
Det är hennes födelsedag i morgon .
Det är hans födelsedag i morgon .
I morgon är det hans födelsedag .
Han har vackra ögon .
Det är dags att åka .
Det är dags att gå .
Om jag var du skulle jag fråga honom .
Om jag var du skulle jag fråga henne .
Om jag vore du skulle jag fråga honom .
Om jag vore du skulle jag fråga henne .
Treviri är Tysklands äldsta stad .
Det var en märklig natt .
Det var en underlig natt .
Han är stolt över att hans son blev läkare .
Hon är stolt över att hennes son blev läkare .
Mary påstod att väskan var en present från hennes man .
Mary påstod att väskan var en gåva från hennes man .
Det var en skänk från ovan .
Ingenting är sant ; allt är tillåtet .
Du har stavat mitt namn fel .
Ni har stavat mitt namn fel .
Du har felstavat mitt namn .
Ni har felstavat mitt namn .
Du har stavat fel på mitt namn .
Ni har stavat fel på mitt namn .
Bussen är tom , och ändå sätter han sig bredvid mig .
Är du hungrig ?
Är ni hungriga ?
Omväxling förnöjer .
Varför är ni på det här skeppet ?
Vill ni inte simma idag ?
Hon går sällan , om någonsin , ensam på bio .
Hon hungrade efter närhet .
Var snäll och avbryt mig inte .
Jag vill inte leka .
Jag vill inte spela .
Vi ska inte på semester .
Ring polisen .
Ring snuten .
Håll utkik efter en skallig och svettig kille .
Gav du dricks ?
Hon är en fanatiker .
Ta reda på vem Tom har pratat med .
Jag får svår prestationsångest före jag ska hålla ett tal .
Vänta , skjut inte !
Jag såg en gammal film på tv .
När jag öppnade dörren hade jag sönder låset .
Tillsätt naturell yoghurt och sojamjölk .
Jag kan springa lika snabbt som Bill .
Jag måste hjälpa honom .
Jag har inga lektioner idag .
Är det något fel på dina ögon ?
Smittar det ?
Jag har ingen kommentar .
Ett slukhål har bildats mitt i motorvägen .
Hur kan folk sova på planet ?
Hur lyckas folk sova på planet ?
Säg mig vad du äter , så ska jag säga dig vad du är .
Jag kan inte läsa franska , inte heller kan jag tala det .
Det här är en läsvärd bok .
Vad står " PTA " för ?
Jag vet att han observerar mig .
Sluta prata om min familj .
Det är det som är kruxet .
Varför är ni på detta skepp ?
Varför är du på detta skepp ?
England och Skottland är grannar .
Du aviseras via e-brev .
Du kan välja att antingen aviseras genom en avi i brevlådan , eller ett sms direkt i din telefon .
Hon sjöng a vista .
Morötter är rika på A-vitamin .
De var tvungna att göra avkall på semesterresan .
Han kastade av sig kläderna direkt innanför dörren .
Ännu en dag är avklarad .
Jag klädde av mig och hoppade in i duschen .
Jag klädde av mig och kröp till kojs .
Var ligger herrarnas avklädningsrum ?
Hon har svårt att koppla av .
Efter en stressig jobbvecka kan det vara svårt att koppla av .
Nu ska jag passa på att koppla av en stund .
De valde att avkorta praktiktiden till tre veckor .
De lastade av bilen och bar upp varorna till lägenheten .
Finska språket har många otroligt produktiva avledningsändelser .
Många av finskans avledningsändelser är mycket mer produktiva än deras svenska motsvarigheter .
Han försökte att avleda uppmärksamheten .
Hennes konstiga beteende var bara en avledningsmanöver .
Han avled förra veckan .
De var tvungna att avliva den svårt sjuka hunden .
Hon spolade ned resterna av innehållet i flaskan i avloppet .
Hon spolade ned resterna av flaskans innehåll i avloppet .
Vi använder endast 10 % av vår hjärna .
Hur löser jag det här problemet ?
Hur löser jag detta problem ?
Hur kan jag lösa det här problemet ?
Hur kan jag lösa detta problem ?
Jag kan inte läsa skrivstil , så kan du vara snäll och texta ?
Hon säljer en ny hatt .
Tom verkar inte komma åt sina data .
Tom verkar inte komma åt sin data .
Du ser ut som en liten flicka i den klänningen .
Jag ska spela fotboll efter skolan .
Tom väntar .
Jag behövde dig .
Jag behövde er .
Hon gick in på sitt rum för att byta klänning .
Hon gick in på sitt rum för att byta kjol .
Janet köpte en klänning och en blus .
Janet köpte en klänning och en skjorta .
Janet köpte en kjol och en blus .
Janet köpte en kjol och en skjorta .
Jag vill köpa den här kjolen .
Jag vill köpa den här klänningen .
Jag har fler kjolar än min storasyster .
Jag har fler klänningar än min storasyster .
Jag tycker inte om ägg .
Jag gillar inte ägg .
Den här röda hatten matchar hennes kjol .
Den här röda hatten matchar hennes klänning .
Den här klänningen passar dig .
Den här kjolen passar dig .
Kavla upp din högerärm .
Jag är upprörd .
Jag önskar att jag kunde simma lika långt som han .
Tom är plastikkirurg .
När pappa kom hem satt jag och tittade på tv .
En katt låg och sov i bastrumman .
Jag vill ha tillbaka mina tjugo dollar .
Vem hatar dig ?
Vilka är det som hatar dig ?
Vem hatar er ?
Vilka är det som hatar er ?
Du kan inte se .
Du får inte se .
Jag är din bror .
Jag är er bror .
Vem förrådde oss ?
Hon vaknade .
Han kanske inte är ung .
Var snäll och spika igen fönstren .
Kom ihåg att följa med mig och fiska på söndag .
Har du någonsin tvättat din bil ?
Har ni någonsin tvättat er bil ?
Vem dog ?
Vem har dött ?
Klockan är sju i London nu .
Hon är sju i London nu .
Han är ett matematiskt geni .
Solen är vit .
John borde vara här när som helst nu .
Försök att inte äta för mycket .
Varför köpte du en blomma ?
De bor i ett nytt hus nära parken .
Kan du hämta mig på stationen ?
Kan ni hämta mig på stationen ?
Du har rätt , Tom .
Kan du kolla om telefonen är trasig ?
Jag fattar inte .
Du fattar inte , eller hur ?
Jag fattar fortfarande inte .
Till min förvåning var han bra på att sjunga .
Han behandlar mig som ett barn .
Du får inte röka .
Två gånger sju är fjorton .
Texas är nästan dubbelt så stort som Japan .
Jag behövde det här .
Det här är brevet från min vän .
Ni fattar inte , eller hur ?
Hur kan jag vara så glömsk ?
Jag glömmer alltid saker till höger och vänster !
Du måste vara Tim Norton .
Pappa är inte hemma .
Seansdeltagare försöker få kontakt med de döda .
Förlåt , jag hade inte med det att göra .
Hon valde ut en rosa skjorta för mig att prova .
Ni får inte röka .
Att bo i en storstad har många fördelar .
Tom försvann .
Adressen på det här paketet är fel .
Jag har en vän vars far är kapten på ett stort skepp .
Hur träffade du honom ?
Du är min enda glädje .
Tom var tokförälskad i Mary .
Han befordrades till överste .
Jag flyttar inte .
Jag flyttar mig inte .
Jag flyttar inte på mig .
De såg förskräckta ut .
Nej , det här pappret är inte vitt .
Vissa kvinnor rakar inte benen .
Vissa kvinnor rakar inte sina ben .
Somliga kvinnor rakar inte benen .
Somliga kvinnor rakar inte sina ben .
Det här är en snuskig film .
Han frågade mig vem jag var .
Hur många ingenjörer deltog i konferensen ?
Du är Toms favorit .
Kan du vara snäll och låsa dörren ?
Kan ni vara snälla och låsa dörren ?
Kan du låsa dörren är du snäll ?
Kan ni låsa dörren är ni snälla ?
De andra barnen kallar henne Piggy .
De andra barnen kallar henne Nasse .
Jane slutade samla på nallar vid tjugo års ålder .
Försvinn från min gräsmatta !
Var inte en sådan surpuppa !
Tom åkte tillbaka .
Tom gick tillbaka .
Vädret ska bli bättre imorgon .
Nästan alla hundar lever .
Jag vill städa huset innan mina föräldrar kommer tillbaka .
Hon bestämde sig för att säga upp sig från sitt jobb .
Vi blev goda vänner .
Vi drack lite vin .
De kommer att göra det .
Magsmärtorna är borta .
Det var intressant .
Hotellet har en hemtrevlig atmosfär .
Kan du höra mig ?
Kan ni höra mig ?
Jag använder det varenda dag .
Hon tittade på några klänningar och valde ut den dyraste .
Vinden blåste hela dagen .
Har du ingenting att göra ?
Har inte du något att göra ?
Har ni ingenting att göra ?
Har inte ni något att göra ?
Det stör mig att hon alltid är sen .
Jag tappade kontrollen .
Hon gjorde så gott hon kunde .
Ring mig senare .
Såg du gårdagens avsnitt ?
Jag hade varit på sjukhuset innan du kom .
Det går inte att förutsäga vad som kommer att hända nästa år .
Han fällde en grötmyndig kommentar .
Markku har hjälpt mig på många sätt .
Att lära sig ett främmande språk kräver stort tålamod .
Jag lär mig tyska .
Är allt där ?
Ung som han är kan han arbeta hela dagen lång .
Ge mig tre kritor .
Våren är kommen .
Ingen rök utan eld .
Och vad ska vi göra nu ?
Och vad gör vi nu ?
Jag håller med Tom .
Vem håller du på ?
Vem hejar du på ?
Vilka håller du på ?
Vilka hejar du på ?
Hon har självmordstankar .
Var är han född och uppvuxen ?
Jag har inget med brottet att göra .
Du måste få tillräckligt med sömn .
Jag ska till Paris .
Hon slog ihjäl honom med en golfklubba .
Jag känner mig sårbar .
Ge henne det här brevet när hon kommer .
Herr Wang kom till Japan för att studera japanska .
Det här är mitt skepp .
Varför följer du efter mig ?
Varför förföljer du mig ?
Varför förföljer ni mig ?
Varför följer ni efter mig ?
Jag köpte en ny handväska .
Vart tog han vägen ?
Vart tog hon vägen ?
Vart tog de vägen ?
Det startade en kedjereaktion .
Vad vill du bli när du blir stor ?
Han skrålade som en hes kråka .
Jag måste gå på min kusins dop .
Hjälp mig bygga färdigt den här sorkstegen så ska jag bjuda dig på middag .
Det går fint !
Han kör utan körkort .
Jag hoppas att det här är början på en vacker vänskap .
Vart gick hon ?
Tom sa att han ville vara här .
Tom sade att han ville vara här .
Han är arton månader gammal .
Min mamma jobbar på fabrik .
Han gick inte upp tidigt .
Han steg inte upp tidigt .
Jag går till skolan på lördag .
Mötet avlystes .
De avlyste mötet .
De visste inte om att de var avlyssnade .
Deras samtal avlyssnades .
Hur ofta lyssnar du av röstbrevlådan ?
Hon fick ett avlångt paket .
Kungafamiljen avlade ett besök på ett av stadens många museer .
Han har avlagt läkarexamen .
Dessa dagar känns sommaren väldigt avlägsen .
Hon ärvde pengar av en avlägsen släkting .
Förövaren avlägsnades från platsen .
Han avläste temperaturen på termometern och skrev upp den i sin loggbok .
I morgon är det avlöningsdag .
Vem ska avlösa henne när hon inte orkar längre ?
Här kommer avlösning .
Hunden kom tillbaka helt avmagrad efter två veckor på rymmen .
Har ni avmaskat valpen ?
Vi befinner oss i en ekonomisk avmattningsperiod .
Den homofobiska retoriken har avmattats med åren .
Nu ska jag avnjuta en kopp te .
Han har en mycket avog hållning till unionen .
Han har en mycket avog inställning till unionen .
Att hitta en perfekt avokado i en mataffär är som att hitta en nål i en höstack .
Tom bad Maria att öppna fönstret .
Det är fruktansvärt dyrt .
Jag har alltid en ordbok nära till hands .
Man stöter på japanska turister överallt .
Han har en vit katt .
Han är amerikan ut i fingerspetsarna .
Hon är tvilling .
Klockan var fem i ett när jag gick till sängs .
Klockan var fem i ett när jag gick och la mig .
Klockan var fem i ett när jag gick och lade mig .
Hon var fem i ett när jag gick till sängs .
Hon var fem i ett när jag gick och la mig .
Hon var fem i ett när jag gick och lade mig .
Den tjocka tjejen äter för mycket sötsaker med mycket socker i .
Den tjocka flickan äter för mycket sötsaker med mycket socker i .
Japaner utbyter gåvor för att uttrycka sina känslor .
Tyskland ligger mitt i Europa .
Han motsatte sig planen .
Jag bor i en lägenhet .
Jag bor i lägenhet .
Det var nästan som en dröm .
Tom är förlovad med Marys lillasyster .
Det är precis som jag förväntade mig .
Jag blir hämtad .
Jag blir upphämtad .
Jag blir uppraggad .
Jag håller på att bli uppraggad .
Tom är trogen Mary .
Två personer kommer in på den här biljetten .
Jag var tvungen att ge upp .
Jag fick ge upp .
Jag fick säga upp mig .
Jag var tvungen att säga upp mig .
Hon dukade av bordet efter middagen .
Det sägs att han är den bästa tennisspelaren .
Den väljaren , Mary Johnson , visade sig vara demokrat .
Ingenting är så enkelt som det verkar .
Inget är så enkelt som det verkar .
Och vad sade de till mig ?
Och vad sa de till mig ?
Och vad berättade de för mig ?
Hur länge måste jag stanna här ?
Bilen körde in i ett skyddsräcke .
Jag är inte det minsta förvånad .
John är här om fem minuter .
Hela familjen hjälpte till med att skörda vetet .
Jag önskar att jag hade ett eget rum .
Jag önskar att jag hade ett rum för mig själv .
England åker ut på straffar igen .
Han håller det hemligt .
Åker han buss till skolan ?
Det här är just den ordbok jag har letat efter .
Tom kommer också till festen .
Du är partisk .
Fisk , tack .
Jag kan inte låta det hända .
De kommer att attackera .
De kommer att anfalla .
Du har inget bra minne .
Jag kunde inte fortsätta ljuga för Tom .
Någon stal mitt pass .
Hon pratar engelska som om det vore hennes modersmål .
Var inte barnslig .
Hur länge har du känt Tom ?
Hur länge har ni känt Tom ?
Publiken såg uttråkad ut .
De köpte det .
De köpte den .
Tom och Mary har varit gifta i tre år .
Jag ville bli astrofysiker en gång i tiden .
Hör du mig bra nu ?
Vi vet ingenting om honom .
Gör inte om det .
Hon talar engelska som om det vore hennes modersmål .
Det är just den här ordboken som jag har letat efter .
Tom är Mary trogen .
Detta kan inte undvikas .
Jag vill inte prata om det just nu .
Jag kunde inte stoppa Tom .
Hej !
God morgon !
Jag är inte din fiende .
Jag är inte er fiende .
Du verkar förvånad .
Ni verkar förvånade .
Du verkar vara förvånad .
Ni verkar vara förvånade .
Förlåt , jag förstår inte vad du säger .
Han är inte längre hemma .
Han är inte hemma ännu .
Ta hand om dig !
Stäng dörren .
Boken är på bordet .
Detta är min dator .
Ni har helt rätt .
Håll tummarna för mig !
Huset tillhör honom .
Hur stavar man ditt efternamn ?
Hur stavar man ert efternamn ?
Liisa kom för sent .
Du är så ondskefull !
Ni är så ondskefulla !
Jag talar klingonska med er .
Jag är en klingonsk krigare .
Han reste sig och gick .
Du ljuger ju bara .
Ni ljuger ju bara .
De togs till fånga .
Hovet städslade en ny städerska .
Var hänsynslös .
Var hänsynslösa .
Använd en skalpell , inte en yxa .
Den där helvilda kackerlackan förfular den så kallade roboten .
Behöver ni hjälp med att bära något ?
Era skor är här .
Ingen kommer att klandra dig .
Ingen kommer att beskylla dig .
Ingen kommer att klandra er .
Ingen kommer att beskylla er .
Tack !
Du är fantastisk !
Tack !
Ni är fantastiska !
Jag kommer inte att följa med dig .
Skynda dig , tåget stannar bara här en kort stund .
Skynda er , tåget stannar bara här en kort stund .
Jag tänker inte lyssna på dig .
Tycker du att jag är larvig ?
Tycker ni att jag är larvig ?
Det här bordet saknar ett hörn .
Detta bord saknar ett hörn .
Alla har kommit nu .
Det är ingen som saknas .
Ingen saknas .
Hinduismen är en polyteistisk religion .
Du är ju helt otrolig !
Du såg lite förströdd ut i dag .
Denna bok är endast för referens .
Utbudet av skor här överstiger efterfrågan .
Efterfesten var i full gång .
Hon vänsterprasslar med grannen .
Hon är otrogen med grannen .
Han talar alltid om gamla barndomsminnen .
Det kan jag inte dra mig till minnes att jag sagt .
Han är väldigt gammalmodig .
Hon är väldigt gammalmodig .
Detta är ett föråldrat tankesätt .
Har du cykelhjälm på dig ?
Brukar du använda cykelhjälm ?
Vi är släkt .
Han är en släkting till mig .
Hon är en släkting till honom .
Du kan äta äpplena med skalet på .
Han drack tre flaskor på raken .
Vi förenas av gemensamma erfarenheter .
Vi utbytte erfarenheter över en kopp kaffe .
Du har ingen aning om vad jag har gått igenom .
Han är utom fara nu .
Det finns en risk för regn i morgon .
Det finns en risk för att han inte kommer .
Skulle du möjligen kunna ha sagt fel ?
Var och en sköter sitt .
Lokalen har nu legat i träda ett tag .
Hon lever ett bekymmerslöst liv .
Jag blev nedkyld av vinden .
Hon somnade så fort hon la sig ner .
Hon somnade så fort som hon lade sig ned .
Bry dig inte om vad andra människor tycker .
Så är det med den saken .
De liknar varandra väldigt mycket .
Han har stukat långfingret .
Det där är skitsnack .
Det där är nonsens .
Kan jag få er uppmärksamhet i två sekunder ?
Sverige är en demokrati .
Sverige är ett folkstyre .
Jag kan följa dig en bit på vägen .
Har du sett vad det blåser ute ?
Vilken stank !
De färdades med båt .
Hon älskar stark mat .
Okej , det går väl för sig den här gången .
Jag har ingen aning om vad han ägnar sig åt nuförtiden .
Jordens öknar breder ut sig .
Gamarna cirkulerade ovanför den stupade antilopen .
Han är noga med vad han tar på sig .
Vi har en del saker att klargöra .
De ska träffas för att göra upp .
Stockholm är Sveriges huvudstad .
Jag är nykter .
Vilken är jordens största öken ?
Vilken är jordens snabbast växande öken ?
Han är klipsk .
Han är snabbtänkt .
Deras framträdande var överlägset .
Till slut fattade de vad vi menade .
Till slut förstod de vad vi menade .
Du har ingenting med detta att göra .
Detta har ingenting med dig att göra .
Hur mår du i dag ?
Känns det bättre nu när du sovit en stund ?
Varför går du inte och lägger dig lite tidigare om kvällarna ?
Denna dator har ett svenskt tangentbord .
Hon har köpt nya hörlurar .
Du måste plugga in kontakten först .
Varför tittar du på mig så konstigt ?
Lagar du middag till mig tills jag kommer hem ?
Hur många gånger ska jag behöva upprepa det här för dig ?
Spelningen var fantastisk rakt igenom .
Hur många tårtbitar åt du ?
Landets ekonomi kollapsade .
Hyllan och alla böcker som stod på den kom ned med ett brak .
Han är en riktig kuf .
Har du något käk ?
Den är ju kruttorr .
Den är ju snustorr .
Den är ju torr som ett fnöske .
Vilken spelevink han är .
Finns det persienner i fönstren ?
Han är aldrig till någon nytta .
I dag har ni varit till stor nytta .
Det är verkligen inte mödan värt .
Det ska snart tryckas upp sedlar med nya motiv .
Något glimmade till i ögonvrån .
Han har ingen ryggrad .
Han är alltid så beskedlig .
Han var inte medgörlig .
Det är viktigt att äta en balanserad kost .
Det står ett spöklikt hus uppe på kullen .
Snön ligger fortfarande på backen .
Snön ligger fortfarande på marken .
Brukar du använda hårsprej ?
Brukar du använda hårspray ?
Hon armbågade sig fram i trängseln .
Det är helt ofattbart .
Det är helt obegripligt .
Han brukar ta färjan mellan Helsingfors och Stockholm .
Gå och kamma dig !
Hur kan ni gräla om en slik sak ?
Han drog en suck av lättnad .
Han släppte sakta upp kopplingen och for iväg .
Den arga hästen sparkade bakut .
Som barn samlade han på skalbaggar .
Detta är ett mycket glesbefolkat område .
De försökte skaka av sig sin förföljare .
Hon avrättades genom hängning .
Nu har datorn hängt sig igen .
Maria studerar socialpsykologi och nu för tiden utforskar hon den europeiska transnationella blogosfärens utveckling .
Han är inte arg .
Vad är det här för skit ?
Han är inte galen .
Varför är hunden här ?
Så synd att ni inte kunde komma .
Skulle du kunna ge oss ett råd ?
Jag vore tacksam för ett snabbt svar och ber dig kontakta mig per mobil .
Några takpannor är spruckna och måste bytas ut .
Mary cyklar på hennes cykel .
Tyvärr hinner jag inte , jag är mycket upptagen just nu .
Jag njuter av min ledighet och bara kopplar av .
När kommer du och hälsa på mig i Sverige ?
Jag ljög för dig .
Jag ljög för er .
Du skrämmer mig inte .
Ni skrämmer mig inte .
Du håller på att bli lat !
Ni håller på att bli lata !
Du är tyst .
Var tyst .
Du ska vara tyst .
Det skickades från min iPhone .
För inte oväsen här .
Hon vet varken hans telefonnummer eller adress .
Du kan gå om du vill .
Ni kan gå om ni vill .
Sover du ?
Jag gör dig nervös , inte sant ?
Jag gör er nervösa , inte sant ?
Jag fick dig att skratta , eller hur ?
Jag fick er att skratta , eller hur ?
Jag fick dig att känna dig obekväm , inte sant ?
Jag har gjort kaffe åt dig .
Jag gjorde kaffe åt dig .
Jag har gjort kaffe åt er .
Jag gjorde kaffe åt er .
Rappakalja pratar jag bäst .
Jag vill inte ha dig här .
Jag vill inte ha er här .
Många av eleverna var trötta .
Jag vet inte om han skulle ha gjort det för mig .
Jag vill veta vad som är roligt .
Jag vill veta vad som är så roligt .
Jag vill veta vad det är som är roligt .
Jag vill veta vad det är som är så roligt .
Tio år har gått sedan jag kom hit .
Det har gått tio år sedan jag kom hit .
Det är galet varmt idag .
Ni är alla bjudna .
Det här är Carrie Underwoods senaste album .
Han hörde illa och kunde inte gå .
Vem har vi att tacka för penicillinets upptäckt ?
Jag sade aldrig att det inte vad en bra idé .
Tom lär sig engelska .
Jag sa aldrig att det inte var en bra idé .
Ingenting spelar egentligen någon roll .
Hade du roligt i helgen ?
Boken kostar fyra dollar .
Hans far vigde sitt liv åt vetenskapen .
Jag vill tillbaka nu .
Matchen kan ha skjutits upp till nästa vecka .
Hon skulle ha gjort det redan .
Hon skulle ha gjort det allaredan .
Han skulle ha gjort det allaredan .
Han skulle ha gjort det redan .
Tom och Mary verkar inte hungriga .
Tom och Mary verkar inte vara hungriga .
De ville inte lyssna .
Ingen gjorde något annat än att dansa .
Jag kan köra .
Engelska är svårt , inte sant ?
Engelska är svårt , eller hur ?
Titta på katten .
Vi åker om en vecka idag .
Kom och träffa några av dina nya klasskamrater .
Jag måste låna lite pengar .
Rökning kan orsaka impotens .
Jag hoppas verkligen att du har rätt .
Jag hoppas verkligen att ni har rätt .
Han vann allt .
Jag minns allt du säger till mig .
Kan du tala esperanto ?
Kan ni tala esperanto ?
Hur fattar du dina beslut ?
Hur fattar ni era beslut ?
Vad ska du med pengarna till ?
Kan ni tala japanska ?
Hon är lika lång som du .
Bladen är gula .
Mannen , som har jackan på sig , är Freddy .
Flickan som heter Inge är från Hamburg .
Det svenska kungahuset har sedan länge enbart representiva och ceremoniella funktioner .
Kollegorna från it-avdelningen är alltid sysselsatta med något annat och har ofta inte tid att ställa upp .
Dessa böcker kan jag rekommendera .
Ett lågtrycksområde täcker hela Skandinavien med växlande vind och molnighet .
Detta är en blyertspenna .
Ormen frestade Eva .
Ibland är det viktigt att fatta ett snabbt beslut .
Jag låtsades arbeta .
Min mor älskar musik .
Du borde fråga honom om råd .
Hon är gift med en tandläkare .
Han är gift med en tandläkare .
Det var alla tiders hur du pratade med henne .
Jag kan inte låta bli att än en gång betona den pedagogiska aspekten av den rapport vi behandlar .
Oj , förlåt !
Jag blandade ihop dig med din syster .
Jag är råkostare .
Detta är ganska dyrt .
Har du en ordbok med dig ?
Det kan jag se med blotta ögat .
Alla hoppades att hon skulle vinna .
Juvelen stals under natten .
Kan du ge mig en filt ?
Jag träffade just henne på gatan .
Mannen åt bröd .
Fader vår , som är i himlen !
Helgat blive ditt namn , komme ditt rike !
Ske din vilja på jorden , liksom den sker i himlen !
Ge oss idag vårt bröd för dagen ; och förlat oss våra skulder , såsom också vi förlåter dem , som står i skuld till oss ; och för oss inte in i frestelse , utan fräls oss från den onde .
Printempo ekvenos .
Jag förstår dig !
Jag förstår er !
En ängslig mor har skarpa ögon .
Jag tackar dig .
Det sägs att Liisa är sjuk .
Jag tackar er .
Har du ätit frukost ?
Har ni ätit frukost ?
Jag vill inte att arbeta under dessa betingelser .
Liisa hade många gånger väntat att Markku skulle säga just dessa ord .
De överraskade henne inte .
Det var tyst mellan dem några minuter .
Markku ville trösta Liisa .
Hur är det med dig ?
Du ser för hemsk ut !
Varför är du så förbannat känslig ?
Nu pratar du fullkomlig smörja .
Vi kommer aldrig överens .
Ting som förr haft betydelse för honom omfattade han med likgiltighet .
Äh , tyst med dig .
Husen brinner .
Mår du inte bra ?
Det är inte billigt .
Jag planerar att tala fler än 20 språk år 2015 .
Jag tycker vi borde göra mer än så .
De fulla sjömännen har ställt till med elände inne i baren .
Jag ställer alarmklockan så att jag inte kommer för sent till jobbet imorgon .
Han flydde från teatern efter mordet .
Herregud , jag kommer komma för sent till lektionen .
Han är helt hopplöst dålig .
Vi är ganska säkra .
Tom beslutade sig för att börja med flugfiske .
Tom är en eldslukare .
Hon kan bara lita på honom .
Vi tappade bort tornet när vi gick in i byn .
Jag gillar att ta mitt block och min penna och åka till kusten för att skissa .
Jag vet inte om vi kan hjälpa dig eller inte .
Bor dem i Algeriet ?
Bränslenivån är under tom.
Sockret är inne i påsen .
Jag tycker inte att hans prestation var något vidare bra .
Ett mynt ramlade ut ur hans ficka .
Kameran som du köpte är bättre än min .
Han är en väldigt hälsosam person .
Han fick malaria medan han bodde i djungeln .
Jag dricker inte champagne .
Jag vill veta exakt vad det är som händer .
Tom blev trött på att alltid behöva betala notan varenda gång han gick ut med Mary .
Hon pratar om Paris som om hon har varit där flera gånger .
Raketen är i omloppsbana runt månen .
Jag gick inte .
Dessa fenomen inträffar , men sällan .
Min far fick mig att tvätta bilen .
Jag vill ha en förklaring .
Tom är en präst .
Jag ville inte spendera mer tid på att arbeta med det där projektet .
Han greps för skattefusk .
Låt oss berätta allt vi vet .
Skadorna från översvämningen räknas bli tio miljoner dollar .
Det vore inte så dumt .
Grattis på födelsedagen .
Jag har ingen flickvän .
Jag är från Brasilien .
Trevligt att träffas .
Han ådrog sig malaria när han bodde i djungeln .
Jag vill inte arbeta under dessa omständigheter .
Jag träffade henne just på gatan .
Jag träffade precis henne på gatan .
Jag träffade henne precis på gatan .
Det här är ganska dyrt .
Det har blivit mycket varmare .
Res dig när ditt namn ropas upp .
Det där är inte billigt .
Raketen ligger i omloppsbana runt månen .
Vi använder endast 10 % av hjärnan .
Vi använder endast tio procent av hjärnan .
Jag vill bara hjälpa er .
Jag vill bara hjälpa dig .
Peter ser väldigt ung ut .
Jag har coola kläder och coola solglasögon på mig .
De olympiska spelen anordnas var fjärde år .
I så fall tror jag att du måste komma i dag .
Alla i bilden ler glatt .
" Tycker du om att resa ? "
" Ja , det gör jag . "
Meddela mig när du slutar .
Du kritiserar alltid mig !
Han åker vanligtvis till skolan med buss .
Hon åker vanligtvis till skolan med buss .
Lejonet rev hundstackaren bokstavligen i stycken .
Jag har ingen lust att gå ut i kväll .
Jag känner inte för att gå ut i kväll .
Skulle ni vilja ha te eller kaffe ?
Det är ett för svårt problem för mig att lösa .
Jag tror att vi glömde någonting .
Jag vill bara vara din vän , ingenting mer .
Är det här franska ?
Är det här franskt ?
Är det här fransk ?
Jag vet att du är rädd för att flyga , men att flyga är inte farligt .
Grannarna var fiender under flera år .
Jag blev upprörd över Liisas beteende .
Barnet är redan döpt .
Markku utnämndes till professor i teologi .
Jag har inga hemligheter för dig .
Jag ringer dig i kväll .
Jag var där ensam i början , men sedan kom Liisa och Liisas nya vän .
Det var trevligt att göra ingenting .
Liisa är en aktiv och energisk ung kvinna .
Jag tycker det är roligt att gå på en promenad .
Jag tycker det är bra att promenera .
Det kan vara .
Han kan inte ha sagt det .
Vilka slutsatser kan dras av detta ?
Det är bisarrt .
Jag tycker att det är roligt att promenera .
Det kan hända .
Det är ju inte så tragiskt .
Nu är jag en riktig gubbe .
Jag blandar mig inte i det .
Använd ditt självförtroende , men aldrig visa upp den för mycket !
Ett av mina barn föddes med någon okänd sjukdom .
Tre av mina barn dog .
Faktiskt kan jag inte riktigt beskriva hur det kändes då .
Det är ganska lätt att tappa tron på att man duger .
Mormor har varit på besök några dagar .
Hur kan man vara så dum ?
Polisen sade att jag måste spärra mitt bankomatkort .
Liisa säger att hon är frisk igen .
Tyvärr kan jag inte komma i kväll .
Markku är en riktigt god vän .
Det smakade bra .
Ett skrattande barn öppnade dörren .
Vad talar du för språk ?
Hur dags äter du frukost ?
Liisa och Markku tycker mycket om varandra .
Flickan som heter Liisa är från Villmanstrand .
Vi hade en lång period av fint väder .
Det är en utmärkt idé !
Jag fick en fantastisk idé .
Jag fick en underbar idé .
Vilka språk talar du ?
Polisen sa att jag måste spärra mitt bankomatkort .
Betty slog ihjäl sin egen mor .
Betty dödade sin egen mor .
Han är en dålig chaufför .
Jag föredrar att gå till fots framför att vänta på nästa buss .
Vad har han gjort ?
Vad har hon gjort ?
Nu är han ombord på skeppet .
Han är inte lång , men stark .
Tom kan köra bil .
Jag förlorade allt jag hade .
Jag förlorade allt som jag hade .
Jag har två barn .
Varje elev har tillgång till biblioteket .
Han har ett hjärta av sten .
Atombomber är en fara för mänskligheten .
Hans hälsa blir sämre och sämre .
Hans hälsa är sämre och sämre .
Jag vet var Tom arbetar .
Jag vet var Tom jobbar .
Jag vet inte vad jag ska göra nu .
Han är rik och mäktig .
Har du två böcker ?
Min bror har fångat en stor fisk .
Det finns en annan möjlighet också .
Jag vet inte vad ni vill att jag ska säga .
Jag vet inte vad du vill att jag ska säga .
Var tolerant .
Var toleranta .
Det hände egentligen inte .
Markku bestämde att han inte skulle stå till tjänst nästa gång och inte någon annan gång heller .
Jag är klarvaken , tankarna snor runt i huvudet som små silverfiskar .
Var ligger hotellet ?
Sluta prata och lyssna .
Jag har en lön på 300.000 yen per månad .
Jag har ont i ögonen .
Jag läser gärna amerikanska romaner .
Korta kjolar är inte på modet längre .
Amerika har olja i överflöd .
Det ligger en bok på bordet .
Tom ringde .
Jag tror att jag har gjort mitt ; det är din tur nu .
Skällde hunden ?
Kort sagt , jag tycker inte om henne .
Hunden har hållit på och skälla .
Oroa dig inte över det !
Sluta med det !
Jag är .
Kan jag kyssa dig ?
Kristus tros ha utfört många underverk .
Det var omöjligt att hitta ett svar .
Det var omöjligt att finna ett svar .
Hon var tvungen att avreagera sig .
Han avreagerade sig på dörren .
Klicka i rutan nedan för att avregistrera dig från våra mejlutskick .
På avresedagen klev de upp redan halv fyra på morgonen .
Hon skrev en artikel i syfte att avromantisera flygvärdinneyrket .
Summan avrundades uppåt .
Kvällen avrundades med en rundtur i trädgården .
Husväggarna hade mjuka , avrundade former .
Försvaret avrustades kraftigt .
Hon avrådde honom från att kritisera ledningen .
Hon gjorde det mot hans avrådan .
Hennes senaste bok avrättades av landets litteraturkritiker .
Han avrättades året därpå .
Han gjorde det i avsaknad av bättre vetande .
Hon hoppade från en klippavsats .
Han ramlade ned från trappavsatsen .
Jag avsåg inte att såra dig .
Denna bok är avsedd för självstudier .
Vad avser tillvägagångssättet har jag inget att invända .
Hon fäster stort avseende vid folks utseende .
Vi gör aldrig avseende på person .
Det här är i alla avseenden en väldigt ogenomtänkt plan .
Bybornas situation är i många avseenden bättre nu än för tio år sedan .
Företaget förlorade avsevärda summor på förra årets omfattande nyanställning .
Han kommer från en avsides by i norra Sverige .
Det var inte min avsikt .
Hon förolämpade honom avsiktligen .
En ansenlig del av befolkningen vill avskaffa monarkin .
De tog avsked och gick skilda vägar .
Han fick avsked på grått papper .
Den stilige mannen räckte henne handen till avsked .
Han avskedades av disciplinära skäl .
De försökte avskeda honom , men han uppfattade inte vinken .
De hittade en avskild strand där de tillbringade dagen .
Det enda som fanns kvar var lite avskrap i botten på kastrullen .
De försökte avskräcka barnen från att leka i skogen genom att berätta historier om vättar och troll .
Han avskyr lukten av surströmming .
Stark avsky mot landets makthavare gav upphov till våldsamma protester .
Skratta inte !
Korsningen där olyckan inträffade ligger här i närheten .
Får jag kyssa dig ?
Jag tycker helt enkelt inte om henne .
Jag tycker helt enkelt inte om honom .
Var köpte du biljetten ?
Sluta vara så nyfiken .
Filmen var avskyvärd .
Han känner sig avskärmad .
Vi öppnade drickan för tre dagar sedan , så den är garanterat avslagen vid det här laget .
Hon kände sig aningens avslagen efter den långa dagen .
Jag är less på honom och hans avslagna idéer .
Det var en avslappnad atmosfär på festen .
Du kan känna dig fullständigt avslappnad i min närvaro .
Efter idrottandet hade de fem minuters avslappning .
Eleverna fick i uppgift att komma på egna avslappningsövningar .
Eleverna fick i uppgift att hitta på egna avslappningsövningar .
De avslutade midsommarfirandet med ett dopp i sjön .
Hon avslutade föreläsningen med att tacka åhörarna .
Skolavslutningen hålls i kyrkan i år .
Skolavslutningen äger rum i skolans gymnastiksal .
På grund av instabil väderlek förflyttar vi skolavslutningen inomhus istället .
Avslutningsvis vill jag tacka alla som kom och lyssnade .
Ansökan avslogs .
Tidningen avslöjade en väl bevarad hemlighet .
Avslöjandet kom som en chock för alla inblandade .
Bara åsynen av mat fyllde henne med en överrumplande avsmak .
De färdades efter en avsmalnande väg .
Polarisarnas avsmältning ökar år efter år .
Hur många avsnitt har du sett nu ?
Vilket avsnitt är du på ?
Hur långt är pilotavsnittet ?
Trots hennes vänliga ton blev hon avsnoppad av den barska busschauffören .
Jag skulle vilja skicka dessa till Japan .
Hon heter Irina .
Nu är det tio minuter till avspark .
Oron avspeglades i hennes ansikte .
Han avspisade henne på ett ytterst snöpligt sätt .
Det är inte blod .
Det är tomatsås .
Din fråga är ologisk .
Jag sitter inte och äter .
Jag håller inte på och äter .
Atmosfären var alltid avspänd när de träffades och umgicks .
Hon är alltid väldigt lugn och avspänd .
Han är en avspänd kille : alltid fötterna på jorden .
De önskar alla en reell avspänning på Koreahalvön .
Hela området är avspärrat på grund av en polisutredning .
Det är förbjudet att vistas innanför avspärrningarna .
Festen var ett avstamp för det kommande samarbetet .
Efter tågolyckan avstannade all järnvägstrafik under tre dagar .
Olika språk har olika regler för avstavning .
Det svenska ordet " bekvämlighet " avstavas " be-kväm-lig-het " .
På väg till Stockholm gjorde de en avstickare till Västerås .
Det finns en avstjälpningsplats tre kilometer norrut .
Hon klev emellan för att avstyra bråket .
Jag tror jag avstår den här gången .
Jag tror jag avstår denna gång .
Han avstod sin plats i kön till en äldre dam .
För henne är avståndet mellan tanke och handling mycket kort .
Partiledaren uttryckte att tydligt avståndstagande från lokalpolitikernas senaste utspel .
Vi vill ha ett kök med gott om avställningsyta .
Detta kök är otroligt svårt att jobba i , då det helt och hållet saknar avställningsyta .
Regnet avtog .
Småtimmarna smög sig på och vinden avtog .
För varje pust avtog vinden mer och mer .
Styrelseordföranden avtackades med blommor och applåder .
Försov dig inte .
Han ville gifta sig omedelbart .
Jag tror det .
Har det kommit några telefonsamtal till mig ?
Markku satte sitt liv på spel för att rädda Liisa .
Låt mig ge dig ett råd .
Liisa hade inte en aning om vad hon skulle göra .
Hans rop på hjälp dränktes i dånet av vågorna .
Och återigen var han hur full som helst .
Såvitt jag vet är det inte så långt .
Vi träffas på kvällen vid bryggan .
Dagens kvinna utsätts för olika påfrestningar .
Hon måste försöka förena både karriär och familjeliv .
Hans karriär inom företaget var över innan den hade börjat .
Smör görs av mjölk .
Välkommen till Wikipedia , den fria encyklopedin som alla kan redigera .
Så vitt jag vet är det inte så långt .
Jag begick ett allvarligt misstag på provet .
Han gick långsamt så att barnet kunde hänga med .
Han gick långsamt så att barnet kunde hinna med .
Han gick sakta så att barnet kunde hinna med .
Han gick sakta så att barnet kunde hänga med .
Han gick sakta så att barnet kunde följa med .
Han misslyckades med att försöka simma över floden .
Jag höll hårt i repet så att jag inte skulle falla .
Många bäckar små gör en stor å .
Har brevbäraren redan kommit ?
Te är en populär dryck över hela världen .
Tom tog någonting .
Jag skulle vilja se dem igen .
Jag skulle vilja träffa dem igen .
Kommer du eller inte ?
Jag stjäl inte .
Varning !
Vått golv .
Vad sägs om en promenad på stranden ?
Vad heter du ?
Är detta en hingst eller ett sto ?
Han odlar många sorters blommor .
Hon odlar många sorters blommor .
Den här genomskinliga vätskan innehåller gift .
Denna genomskinliga vätska innehåller gift .
Det internationella språket interlingue offentliggjordes 1922 under namnet Occidental .
Ring dem i kväll .
Min hund åt min läxa .
Jag tänker , alltså är jag .
Min kniv är vass .
Jag var lärare .
Det är ingen hemlighet .
Mitt glas är fullt .
Det var aldrig svårt för oss att hitta något att prata om .
Hon kunde inte sluta le .
Varför slutar du inte ?
Varför slutar ni inte ?
Är det moraliskt fel att äta kött ?
Tom undrar om det är sant .
Han kanske ljög för mig .
Hon kanske ljög för mig .
Jag är seriös .
Kan jag komma ut ?
Jag måste gå nu .
Hon var i ett kritiskt tillstånd .
Vi ses !
På återseende !
Vi håller kontakt .
Han bor i det där huset .
Hon bor i det där huset .
Han bor i huset där borta .
Hon bor i huset där borta .
Varför har du inte klänning på dig ?
Ta på dig en klänning då .
Han ramade in fotografiet och hängde upp det ovanför sängen .
Hon gav henne ett kvitto som hon hade skrivit sitt telefonnummer på .
Från den här vinkeln ser jag inte ens halva duken .
Du glömde din mobilladdare hos oss i går .
Skicka den på posten så får jag den om en dag eller två .
Någon måste ha tagit mitt paraply av misstag .
På tal om herr Tanaka , har du sett honom på sistone ?
Jimmy insisterade på att jag skulle ta honom till zoot .
Mitt hus ligger i norra delen av staden .
Min pappa insisterade på att vi skulle vänta på tåget .
Min far insisterade på att vi skulle vänta på tåget .
Skulle du kunna förklara reglerna för mig , tack ?
Skulle ni kunna förklara reglerna för mig , tack ?
De skyndade sig till olycksplatsen .
Båda mina systrar är gifta .
Du måste inte komma hit varje dag .
Ni måste inte komma hit varje dag .
Han är konstig ibland .
Vi uppfattar inte saker som dom är , utan som vi är .
Frågan är inte vad jag kan vinna utan vad jag har att förlora .
Hon pratar inte bara flytande engelska utan också flytande franska .
Han var så upptagen att han skickade sin son istället för att gå själv .
Det viktiga är inte hur en man dör , utan hur han lever .
Framtiden tillhör inte de ängsliga , den tillhör de modiga .
Det är inte en fru jag vill ha , utan en knullkompis .
Vi spelade schack inte så mycket för att vi gillade att spela som för att bara slå ihjäl tiden .
Krig startar inte bara som vintern startar , utan snarare är det människor som startar ett krig .
Hon är inte sjuksköterska , utan läkare .
Ingendera är vacker .
Jag vill bara vara med dig .
Hon var på humör för en promenad .
Varför hände det här ?
Det fanns ingen kvar utom mig .
Jag utgick ifrån att du skulle närvara på mötet .
Han kan mycket väl ha rätt .
Han kan ha rätt .
Där är vackra blommor här och där i trädgården .
Vi iakttog honom tills han var utom synhåll .
Varför vill du att världen ska känna till japanska trädgårdar ?
Kunde du ta det här , tack ?
Toms bil är lätt igenkännbar eftersom det är en stor buckla i den främre stötfångaren .
Jag gillar verkligen hårdkokta ägg .
Han förklädde sig till en kvinna .
En del av uppsatserna är mycket intressanta .
Vi flyttade våra väskor för att ge plats för den gamla damen att sitta ner .
Det finns många städer i det här landet .
Det finns många arter av fiskmås som varierar i storlek .
Det låter som om du är upptagen .
Tom lurade dig .
Har du grävt upp potatisar ?
Jag kommer inte på någonting .
Hon ville veta om fotografen kunde ta bort hatten från bilden .
Jag förlorade henne ur sikte i folksamlingen .
Alkohol löser inga problem .
Vi kan inte prata nu .
Ölglaset är nästan större än dig .
Jag rådde honom att komma tillbaka omedelbart .
Ken läste när jag kom hem .
Jag har en överraskning för dig .
Självklart tycker jag om det .
Vad dom säger är sant .
Det är ett gammalt manuskript .
Hon talar tillräckligt tydligt för att vara lätt att förstå .
Hans systrar så väl som han själv bor nu i Kyoto .
Doktorn sa till herr Smith att sluta röka .
Det är en oklar historia .
Tom ville inte berätta för Mary att han hade förlorat alla hennes pengar .
Det är likartat .
Tom lever ur hand i mun .
Tom visste inte vad han skulle göra härnäst .
Terrorism är den viktigaste faktorn för delningen av ett land och skapandet av självständiga regioner .
Kan du skicka saltet ?
Jag vill hålla mitt rum så prydligt som möjligt .
Han visste inte vad han skulle göra .
Hisaos ansikte var likblekt .
Hon var på vippen att gråta .
Hur lång tid tar det att ta sig till Wien till fots ?
Jag kan göra det härifrån .
Man bör läsa många böcker när man är ung .
Jag letar efter något att tvätta mattan med .
Ser du porträttet ?
Att ta genvägar sparar pengar på kort sikt men förlorar kunder på lång sikt .
Du är avskedad !
Vad undersöker en sovjetolog ?
Vad studerar en sovjetolog ?
Han är en sångare .
Hon är en sångerska .
Det här bordet är vitt .
Den här pennan är bäst .
Det här är inte fisk .
Han vill spela fotboll i eftermiddag .
Det här är en penna .
Vi ser inte saker som de är , utan som vi är .
Hon var gråtfärdig .
Hon var gråtfärdig .
Det är liknande .
Jag har en överraskning åt dig .
Det är likt .
Jag har en överraskning åt er .
Den är liknande .
Den är lik .
Vi ser inte saker som de är , utan som vi är .
Är han här snart ?
Det var det .
Det om det .
Abonnenten du försöker nå kan inte ta ditt samtal just nu .
Vänligen försök igen senare .
Dom bär dyrbara ringar .
Jag har korrigerat misstaget .
Klockan var nästan 2 : 30 när Tom till slut kom hem .
Jag vet att du är arg .
Det kommer aldrig att hända .
Tom låtsades inte veta vart han skulle gå .
De bär dyrbara ringar .
De bär dyra ringar .
Jag brände pappret .
Ingången till toaletten är mycket smutsig .
Åt du något ?
Jag brände papperet .
Hur många gånger ska jag måsta säga det till dig ?
Hur många gånger måste jag säga det till dig ?
Jag är inte läkare .
Ingen skall överleva .
Hur länge tänker du stanna här i Brasilien ?
Du sover i mitt rum .
Jag återvände från skolan .
Jag drack kaffet .
Jag öppnar en låda .
Jag kan inte förstå .
Det här är en bild av min syster .
Emily skriver ett brev .
Bilen är blå .
Jag sjunger en skön sång .
Jag sjunger en sång .
Du kommer att förstå att jag berättar sanningen .
Jag drack inte vattnet .
Emily frågade en fråga .
Europa är en kontinent .
Jag skall gå till stranden .
Det där är ett hjärta .
Mitt hjärta blöder .
Jag skall gå till parken .
Jag har blå ögon .
Jag har röda ögon .
Hassan gick till skolan .
Katten är under bordet .
Han åt äpplet .
Jag skall läsa boken .
Vetenskapen är viktig för våra liv .
Jag tror inte att två språk är tillräckligt .
Jag vill leva i staden .
Jag ser huset .
Hur gammal är din son ?
Hur kan jag få dig att ändra dig ?
Jag måste göra min läxa .
Du måste göra din läxa .
Jag äter en bok .
Jag ska läsa boken .
Jag ska gå till parken .
Är jag fadern ?
Jag ska gå till stranden .
Vi älskar dig så mycket .
Min hund skäller hela tiden .
Jag sjunger en vacker sång .
Det finns ett brev för dig .
Ingen kommer att överleva .
Det nya huset ligger här .
Hon kan simma .
Han kan simma .
Det finns en katt i lådan .
Jag frågar henne en fråga .
Det här är mitt hus .
Jag kan äta .
Jag kan inte äta .
Jag lokaliserar programvaran .
Jag har ett hjärta .
Jag har en katt .
Den här dörren går inte att låsa .
Denna dörr går inte att låsa .
Jag gick inte till skolan .
Den här dörren är inte låsbar .
Denna dörr är inte låsbar .
Jag skall äta äpplet .
Kärleken är en viktig sak .
Jag ska äta äpplet .
Vilket högt nummer !
Jag bor i Qatar .
Det här är en hönsfågel .
Min penna är i min hand .
Jag går och lägger mig klockan tio .
Jag går till jobbet klockan sju .
Ditt blod är rött .
Jag skrev inte ett brev .
Jag går och lägger mig klockan tio .
Emily kan simma .
Jag köpte henne en vacker klänning .
Det här är en liten bok .
Vi vann tävlingen !
Jag förstår dina ord .
Har du en ordbok ?
Jag behöver en bättre ordbok .
Jag vill lära mig svenska .
Jag återvände till huset .
Vill du ha fisk ?
Talar du arabiska ?
Jag talar arabiska .
Han återvänder till sitt hem .
Jag är studerande .
Det här äpplet är rödare .
Jag kommer från Turkiet .
Det ligger en apelsin på bordet .
Det är bäst att du åker hem så snart som möjligt .
Jag tar snart kontakt med dig .
Jag tar kontakt med dig snart .
Åk vart du vill .
Gå vart du vill .
Har du svårt med att förstå vad kvinnor och barn säger till dig ?
Jag vill inte höra några ursäkter .
Vad är din blodgrupp ?
Jag kan leva utan vatten .
Skulle du kunna ögna igenom de där pappren lite ?
Skulle du kunna ögna igenom de där papperen lite ?
Vi hade ingenstans att bo .
Mjölken surnade .
Han verkar aldrig åldras .
Stockholm är Sveriges huvudstad .
Sveriges huvudstad är Stockholm .
Han tror inte att jag förstår hans taktik .
Förresten , var bor du ?
Var bor du , förresten ?
Var bor du nuförtiden ?
Var bor du nu ?
Var är ditt hus ?
Hon är så stor !
Det lyster honom att se de små leka i vattenbrynet .
Vet du hur hon mår ?
Var är de vackraste meningarna ?
Min GPS-navigator fungerar inte utomlands .
Hon grät sig till sömns .
Hon somnade gråtandes .
Hon tog emot sedeln utan att säga någonting .
Katten sover på bordet .
Vilken skola är bäst ?
Jag gick till sjukhuset .
Det finns lite grädde i kylskåpet .
Med vänling hälsning , Silja
Du förtjänar mer .
Du vill ha dom här grejerna , inte sant ?
Han var synligt nervös .
Konferensen kommer att hållas i Tokyo .
Jag var tvungen att hämta någonting från mitt rum .
Jag tror att jag kommer att kunna träffa dig snart .
Hon är fortfarande minderårig .
Han har precis kommit hem .
Det ska bli kallare och snöa senare idag .
Du vill ha de här grejerna , inte sant ?
Har du svårt att gå ner i vikt ?
Brevet är skrivet av flickan .
Någon stal mitt körkort .
Vem är jag ?
Var kommer jag från ?
Finns det liv efter döden ?
Vad är meningen med livet på jorden ?
Låt oss spela volleyboll .
Det finns så många självrättfärdiga människor .
Öga för öga , tand för tand .
Det finns ett fel i meningen .
Jag hörde åskdundret , men såg inte blixten .
Låt oss spatsera litet på stranden .
Detta fält är inte väl odlat .
Jag delar inte din åsikt .
Jag är rädd för höjder .
La Lia Rumantscha är paraplyorganisationen för alla rätoromanska kvinnor och män .
Den vill på ett hållbart sätt främja det rätoromanska språket och dess kultur .
Jag är höjdrädd .
Hon öppnade dörren .
Vi behöver köpa vinäger .
Jag ber om ursäkt för det .
Läraren öppnade lådan och tog ut en boll .
Staden ligger vid havsstranden .
Titta inte på kameran .
De har läst en intressant bok .
Jag kom hem sent .
De lät mig välja en present .
Jag vill se gatorna .
Det var en stor en .
Han blev polis .
Tom bad mig om hjälp .
Varför bryr hon sig inte om mig längre ?
Frukosten serveras klockan sju .
Finns det någon som kan svara ?
Men det är inte det sista tåget , eller ?
Tom kan inte bestämma sig för vilken kamera han ska köpa .
Det finns få webbsidor på tatariska på internet .
Jag vill inte dö !
Grattis !
Detta skickat från min iPhone .
" Du , min herre , är en imperialist ! "
" Och du , min herre , är ett troll ! "
Det starka ljuset störde Markku .
Boken intresserar mig .
Såvitt jag vet är detta inte fallet .
Tom tände bordslampan .
Jag har bra dagar och dåliga dagar .
Mark tog sina saker och gick .
Sanningen att säga , led änkan av magcancer .
Råttan är en gnagare .
Rapporten ansågs vara falsk .
Så vitt jag vet är detta inte fallet .
Är det någon som kan svara ?
Vi har en hel del att prata om .
Markku tillbringar mycket tid framför tv : n .
Jag tror att Tom och John är enäggstvillingar .
Jag kan faktiskt inte svaret .
Jag vet faktiskt inte svaret .
Engelska är , som du vet , i högsta grad ett levande språk .
Engelska är , som ni vet , i högsta grad ett levande språk .
Vi bakar kakor .
Jag fastnade .
De älskade det .
De älskade den .
Hennes ledighetsansökan avslogs .
Jag funderade på planen .
Deras kontrakt går ut i slutet av den här månaden .
Deras kontrakt löper ut i slutet av den här månaden .
Deras kontrakt går ut i slutet på den här månaden .
Deras kontrakt löper ut i slutet på den här månaden .
Han är lika lång som min far .
Han är en av Spaniens mest kända författare .
Hon är orolig för sin vikt .
Hon oroar sig för sin vikt .
Tittar de på oss ?
Jag måste ha passerat stationen medan jag tog en tupplur .
Min mor tar en tupplur varje eftermiddag .
Skynda dig , annars missar du tåget .
Tom är min brorson .
Tom är min systerson .
Jag tycker om att simma , men inte här .
Mitt huvudämne på universitetet var kemi .
Ska vi beställa ?
Hyddan stacks i brand .
Kojan stacks i brand .
Skjulet stacks i brand .
Han stack sitt hus i brand .
Han satte eld på sitt hus .
Mannen satte eld på sig själv .
Han tillverkade en liten hundkoja .
Jag satte upp en liten koja i trädgården .
Kan jag få en kudde ?
Jag behöver en extra kudde .
Den rosa kudden är ren .
Den där dunkudden ser dyr ut .
Min kudde är så mjuk !
Hon kvävde honom med en kudde .
Tom bad om en filt och en kudde .
Tom och Mary hade kuddkrig .
Vilken skitstövel !
Det var oförlåtligt .
Jag börjar tappa tålamodet .
Han gick ut en runda med hunden .
Det var brännbollsturnering på allmänningen .
Nu har jag snart ätit upp , men någon groda har jag då inte sett röken av .
Får jag raka av dina polisonger ?
Var god fyll i enkäten och skicka in den till oss .
Först visste jag inte vad jag skulle göra .
Först visste jag inte vad jag skulle ta mig till .
Hans frånvaro igår berodde på hans förkylning .
Man måste göra vägen lång för att spara tid .
Räven byter pälsen men inte lasterna .
Äta kan man allt man har , men inte berätta allt man vet .
Den som sjunger om somrarna , arbetar om vintrarna .
Folk och väder måste man ta som de är .
Människor utan humor är som ängar utan blommor .
Man blir inte mästare på en dag .
Bra och fort går sällan ihop .
Ett fruktansvärt kaos härskar i vardagsrummet .
Det är läggdags .
Jag vet inte riktigt än .
Jag ska till Paris i helgen .
Vi översatte rapporten från engelska till afrikaans .
Jag gillar österrikisk musik .
Jag tycker om österrikisk musik .
Jag såg Tom för mindre än en timme sen .
Jag såg Tom för mindre än en timme sedan .
Edward Sapir var en amerikansk lingvist .
Han bestämde sig inte för att bli författare förrän han var trettio .
Jag ska prata med Tom när han kommer hem .
Han tog sig friheten att skriva till damen .
Kan du ta hand om våra husdjur medan vi är borta ?
Kan ni ta hand om våra husdjur medan vi är borta ?
Vad gjorde Tom med pengarna ?
Vad gjorde Tom av pengarna ?
Jack då ?
Du då ?
Vill du också ha apelsinjuice ?
Du då ?
Vill du också ha apelsinjos ?
Du då , litar du på den här mannen ?
Ni då , litar ni på den här mannen ?
Du förtjänar det här .
Tom kör .
Vilken tid passar dig ?
Vilken tid passar er ?
Vann du ?
Vann ni ?
Vi lärde oss ryska istället för franska .
Så du ska ingenstans imorgon ?
Jag har många samtal att ringa .
Jag har många beslut att fatta .
Jag vill verkligen tala om för damen som klipper mitt hår att jag inte tycker om att ha lugg .
Han rusade in i rummet .
På två drag kommer Kasparov att ställa motståndaren i schack .
Du har blivit tjock .
Jag försöker komma på varför någon skulle göra något sådant .
Jag försöker komma på varför någon skulle göra någonting sådant .
Jag försöker komma på varför någon skulle få för sig att göra något sådant .
Jag försöker komma på varför någon skulle få för sig att göra någonting sådant .
Vi kan inte hålla med dig på denna punkt .
Jag håller inte med .
Hon är stolt över sin dotter .
Jag är idel öra .
Jag vill inte lägga mig i .
Och det är det !
Han är elva år gammal .
Jag har ett dåligt samvete .
Jag kommer inte ihåg texten .
Jag kommer inte ihåg orden .
Jag minns inte texten .
Jag minns inte orden .
Den här filmen är ett mästerverk .
Rökning är förbjudet .
Hur många kvadrater kan du se ?
Jag har fått en bil .
Detta är första gången som jag är gravid .
Han bodde i Azerbajdzjan i 4 år .
Han är sällan hemma .
Då ska jag se vad jag kan göra !
Kor äter gräs .
Tom är en ganska envis .
Fastighetsmäklaren ljög för paret .
Vi har inte hittat Tom .
Påven Francis återvänder till Rio år 2016 .
Om ni sticker oss , blöda vi icke ?
Du är bara nervös .
Varje morgon läser jag om vädret i tidningen .
Var snäll och kom och hjälp mig .
Jag vill ha en öl .
Mina vänner stod vid min sida under rättegången .
Han kommer aldrig att erkänna sin skuld .
Han kommer aldrig att erkänna att det är hans fel .
Mina vänner svek mig inte under rättegången .
Tom borde definitivt ha fått dödsstraff .
Jag kan inte minnas att jag har bett om din hjälp .
Han dog innan ambulansen kom .
Han stängde dörren .
En nyfödd baby är benägen att bli sjuk .
Hördu , jag vill inte förlora mitt jobb .
Medicinen gjorde underverk för hans hälsa .
Vem arbetar du för ?
Tom är en man med många talanger .
Tom älskar Mary .
Jag njöt av den vackra våren .
För ett ögonblick trodde jag att han hade blivit galen .
Det var nära !
Vad fick dig att komma hit ?
Jag kan inte stå ut med sin fräckhet .
Jag försökte att inte gråta .
Verkligen ?
Om jag bara hade bett om ditt råd .
Jag är inte din fru längre .
Din fru är Tatoeba !
När jag jobbar , dricker jag en massa kaffe .
Man tjänar inte på det i längden .
Du tjänar inte på det i längden .
Liisa kom för tidigt .
Du måste vara försiktig .
Han kommer att vara ledig imorgon .
Tom släckte lampan på nattduksbordet .
Ögonen är själens spegel .
Han är en sefardisk jude .
Jag ska vila mig lite .
Hon var en av de första svenska kvinnor som avlade doktorsexamen i matematik .
Han doktorerade på en avhandling om medeltida kyrkokonst i Norden .
Beslutet överklagades senare till länsstyrelsen .
Jag skulle vilja skicka ett rekommenderat brev .
De genomförde flera studieresor i Norden .
Han etablerade sig snabbt som en av landets mest lästa författare .
Universitetets huvudbyggnad ritades av en ung dansk arkitekt .
Hennes familj flyttade runt en hel del .
Han dömdes till livstids fängelse .
Hon ville avsäga sig sitt amerikanska medborgarskap .
Jag skulle vilja ha en gaffel .
Jag har många språkböcker .
Tom bröt mot reglerna .
Jag skulle vilja skicka ett rek .
Han är ledig i morgon .
Hon är ledig i morgon .
Om du vill köpa ett koppel , gå till en zooaffär .
Jag vill vara ett barn .
Har ni sett den här ?
Vampyren suger mitt blod .
Krig är helvetet .
Jag arbetade .
Jag kan inte bullra .
Barnet sover .
Republikanerna var rasande .
Bron var byggd av romarna .
Du blir tvungen att laga mer mat .
Vem gick du med ?
Enligt tidningen ska det snöa imorgon .
Ingen vill ha ett krig .
Det var ett oförlåtligt misstag .
Kardborre är en tvåårig medicinalväxt .
Hon ljög .
Alla djur är lika .
Varför kan Tom inte komma ?
Vad är grafen ?
Grafen är ett ämne som består av rent kol .
Grafen är 200 gånger starkare än stål .
Huvudstaden i Ukraina är Kiev .
Det är den bästa vi har .
Hon bad sin lärare om råd .
Du måste lyckas där dom största hjältarna har misslyckats .
Fången befanns skyldig .
Tom och Mary var dom två sista att ge sig av .
En del människor tjänar stora pengar ur tomma luften på finansiella transaktioner .
Varför kan vi inte helt enkelt bestämma att alla är stormrika från början ?
Solen lyser även på natten .
Hösten hade kommit till landet .
Pennan är kanske mäktigare än svärdet , men den är då inte mäktigare än pennvässaren .
Var snäll och översätt den här meningen till valfritt språk .
Nadir är när solen står på rakt motsatt sida av jorden .
Det är motsatsen till zenit .
Det Tatoeba framförallt lär en är att man inte ens kan tala sitt modersmål .
Piloten lyckades genomföra en perfekt landning .
Katter finns i många olika storlekar .
President Grant har inte gjort något olaglig .
Han är mycket förstående .
Hon kommer kanske imorgon .
Den här boken är unik på många sätt .
Kung George tog kontroll över kolonin 1752 .
Stationen är två engelska mil bort .
Låt oss stoppa här .
Tom visste inte vad det var meningen att han skulle göra .
Eftersom han är gift , måste han tänka på framtiden .
Den finansiella situationen förvärras vecka för vecka .
Dom här skorna är dyra , och dessutom är dom för små .
Han går vanligtvis hem klockan fem .
Min far lyssnar på klassisk musik .
Jag har en vit katt .
Heather tror mig .
Tom klarar sig jättebra .
Förlåt honom om du kan .
Han är oskyldig .
Tom klarar sig mycket bra .
Produktionen har börjat avta .
Vi börjar mötet när Bob kommer .
Den här pingvinungen är så söt !
Jag föddes med tolv fingrar .
Du måste arbeta snabbt .
Ni måste arbeta snabbt .
Jag ska inte förråda Tom .
Den här byggnaden ska byggas i staden .
Jag vill inte leva med dig .
Jag spelar i trädgården .
Det är inte möjligt .
Spinoza var en panteist .
Lejonet är kungen av djungeln .
En spegel reflekterar ljus .
Jag vill gifta mig med Heather .
Jag föddes och växte upp i landet .
Tom ser verkligen ledsen ut .
Det varierar en hel del .
De allierade kontrollerade alla större irakiska städer .
Vilken lägenhet som helst duger så länge hyran är rimlig .
Jag sköt upp hushållsarbetet några timmar .
Jag sköt upp mitt hushållsarbete några timmar .
Jag sköt på mitt hushållsarbete några timmar .
En bok är tunn och den andra är tjock ; den tjocka har cirka 200 sidor .
Vet du om han kommer till festen ?
Jag får inte gå härifrån .
Jag gick upp för en timme sen .
Vem som än använder den här tandborsten är inte min mor .
Herr Wilson tvingade oss att upprepa meningen flera gånger .
Bar båda hjälmar ?
Snälla ge mig någonting att äta .
Mödrar brukade säga till sina söner att om dom masturberade skulle dom bli blinda .
Klippan är nästan vertikal .
Låt oss hålla kontakten med varandra .
Han arbetar fortfarande i arbetsrummet .
Var täckte du över dom ?
Tom kunde inte besvara en endaste fråga på gårdagens test .
En mans ansikte är hans självbiografi .
En kvinnas ansikte är hennes skönlitterära verk .
Det slog honom aldrig att hon skulle bli arg .
Han är bra på rugby .
Jag har hållit på att skriva det här manuskriptet i ett år .
Han begick många synder i sin ungdom .
Jag lät mina känslor fördunkla mitt omdöme .
Talar Tom flytande franska ?
Jag är trött eftersom jag arbetade för mycket .
Jag lyssnar nästan aldrig på radio .
Jag ska berätta sanningen .
Låt oss tala engelska .
Jag mindes alla .
Tycker du om det ?
Tom moppar golvet .
Den svarta kattungen hoppade för att undvika pölen , och passerade under den angränsande häcken .
Det var hans bil , inte min , som gick sönder igår .
Håll mig informerad tack .
Jag vill inte se dum ut .
Ingen är rik i mitt land .
Jag vill inte verka dum .
Tankar uttrycks genom ord .
Vill du ha mer kakor ?
Fast han är mycket fattig , är han ändå för god för att ljuga .
Du måste kämpa mot den tendensen hos dig .
Tankar uttrycks med hjälp av ord .
Han har ett stort ego .
Knivspetsen är vass .
Jag är i princip lika kvalificerad som Tom .
Han är av naturen en vänlig person och populär hos barnen i området .
Han brände hål i rocken .
Tom kommer inte att göra det .
Om du får någon tid över , använd den och gör dina läxor .
Det beror på , förstår du , att jag har vetat sen länge att han inte är den sortens människa .
Varför är dom rädda ?
Alla rören frös förra vintern .
Den här motorn ger ibland upp andan .
Hon slöt sina ögon .
Har du någonsin sett Buckingham Palace ?
När kommenterade du en mening senast ?
Detta är ett historiskt ögonblick .
Det dom sökte var en man som han själv .
Det är utpressning .
Vad betyder SSSR ?
Jag ville att Tom skulle känna sig som hemma .
Tom såg Mary på TV .
Tom arbetade deltid .
Tom kan inte läsa utan glasögon .
Vem sitter vanligtvis på åsnebänken ?
Detta är intressanta nyheter .
Filmen börjar klockan tio .
Mary är nu en glad liten flicka .
Deras favoritämne var eskatologi .
Att oroa sig är som en gungstol ; det ger en någonting att göra men leder ingenstans .
Om jag då hade kunnat tala franska , hade jag inte fått några problem .
När jag springer , blir jag svettig .
Han är min dubbelgångare .
Hon vill arbeta på ett sjukhus .
Jag talar om dina åtgärder .
Kan jag hjälpa dig ?
Det är förnedrande för henne .
Det kan du vara säker på .
Jag ska aldrig glömma Toms ansikte .
Tom kunde inte öppna dörren .
Afrika är mänsklighetens vagga .
För ögonblicket har vi större problem .
Just nu , har vi större problem .
Vi hade våra skäl .
Du behövs inte .
Ni behövs inte .
Du är överflödig .
Tom minns inte var .
Om du vill , så ring mig på eftermiddagen .
Det är inte för att hon är vacker som jag gillar henne .
Vi genomförde vår utredning med största noggrannhet .
Åh , ta god tid på dig .
Jag har ingen brådska .
Koppen är sprucken .
Vi har inget behov av assistans .
Tom har studerat franska i ungefär tre år .
Inatt var det väldigt varmt och kvavt och jag sov inget vidare .
Tom och Mary var på Johns begravning .
Hon rådde honom att prata om sitt liv i Förenta Staterna .
Toms far är en berömd konstnär .
Jag förmodar att han kommer .
Jag ångrar att jag var så lat under min skoltid .
Det finns ingenting jag kan göra .
" Kunde du hämta en kopp kaffe åt mig ? "
" Visst .
Så gärna . "
Du kan köpa frimärken på vilket postkontor som helst .
Ni kan köpa frimärken på vilket postkontor som helst .
Man kan köpa frimärken på vilket postkontor som helst .
Jag känner henne inte .
Jag vill inte att det ska finnas några lögner mellan oss .
Jag vet inte när han kommer , men när han gör det , kommer han att göra sitt bästa .
Det har gått tre år sedan vi gifte oss .
Tom kunde inte bestämma sig omedelbart .
Han förnekade sin inblandning i historien .
Jag kanske går ut om det slutar regna .
Ut allesammans !
Han är något av en musiker .
Jag tycker att vi borde vänta .
Jag har inte sovit något vidare .
Fråga mig någonting enklare .
Han har en stor restaurang nära sjön .
Det var hans beslut .
Hur många delfiner finns det på detta oceanarium ?
Du kan lika gärna börja omedelbart .
Bergets övre del är snötäckt .
Jag var inte medveten om att Tom hade gjort det .
Huset är mycket gammalt .
Det behöver repareras innan du säljer det .
Huset är mycket gammalt .
Det behöver repareras innan ni säljer det .
Tom talade till Mary från den andra sidan .
Jag är en vegetarian som äter massor av kött .
Hon måste vara död .
Han har inga vänner .
Det är dumt att läsa en sådan tidskrift .
Hon hatade vanilj .
Under den stalinistiska eran blev fångar i koncentrationsläger slavar i statens tjänst .
Robin är Batmans vän .
Jag översätter inte romaner längre .
Håll bollen i rullning .
Jag är emot det .
Jag växte upp i en fattig familj .
Jag visade dem hur man gör det .
Jag talar om ditt handlande .
Jag talar om ditt agerande .
De här skorna är dyra , och dessutom är de för små .
Vi stannar här .
Bron byggdes av romarna .
Snälla sluta !
Jag vill inte att någon ska bli skadad .
Vi är båda galna .
Jag sa att det var ok .
Du kom in i mitt rum .
Ni kom in i mitt rum .
Jag blev nästan påkörd av en bil .
Ingen människa bor i byggnaden .
Ingen man bor i byggnaden .
Vi väntade på båten i många timmar .
Dom var utmärkta .
Det är otroligt .
Han har en bil som jag gav honom .
Det är dags att vi söker nya utmaningar .
Jag är smickrad .
Är vi inte vänner ?
Han sov i bilen .
Tror du att det kommer att regna idag ?
Tror ni att det kommer att regna idag ?
Vad tror du hände här ?
Vad tror ni hände här ?
Du kan inte ersätta kommat med en punkt i den här meningen .
Jag försökte att inte skratta .
Liisa uppförde sig som om hon visste allt .
Jag måste vara försiktig .
Jag ser fram emot det .
Du kan inte döda dig själv genom att hålla andan .
Jag vill tala engelska .
Min engelska är inte god .
Det är felaktigt .
Emily vill arbeta i ett stort företag .
Emily är en gottegris .
Jag talar tyska .
Älskar du henne ?
Hon hade gått till skolan .
Jag kan älska det .
Jag har lärt mig något från den här boken .
Hur kan speglar vara sanna om våra ögon inte är äkta ?
Jag har aldrig röstat .
Jag träffade henne på vägen till skolan .
Han studerar astronomi , eller stjärnlära .
De är korta och smala .
Hon kopierade en mening .
Hon behöver hjälp .
Hon vattnade ett träd .
Hon vann en telefon .
Hon bar en mask .
Hon skrev en kort berättelse .
Hon tvättade en matta .
Hon översatte en dikt .
Hur mår du , Mike ?
Ursäkta mig , jag har en förfrågan .
Vi hyrde en lägenhet .
Livet är som en stor huvudväg .
Kvinnan äter bröd .
Jag läser den här tidningen .
Det finns en pojke i det här rummet .
Det finns en hund i det här rummet .
Jag skulle vilja köpa en hund .
Jag kramade Emily .
Emily kramade mig .
Jag ska berätta det för Emily .
Emily ska berätta det för Melanie .
Emily skrev meningen .
Jag åkte till Danmark .
Jag åkte till Sverige .
Jag åkte till Norge .
Vi gick till stranden .
Hon sjöng en sång .
Med till visshet gränsande sannolikhet hade mannen begått självmord .
Markku ville inte ligga sin far till last .
Oroa dig inte för mig .
Liisa var allmänt omtyckt och hade lätt för att skratta och skämta .
Liisa stirrade förbluffat på Markku .
Det fanns inte mer att säga om saken .
Du är här för att sköta ditt jobb .
Markku rynkade ögonbrynen .
Jag har inte den blekaste aning .
Jag har nu blivit döden , världarnas förintare .
Markku rynkade på ögonbrynen .
Min engelska är inte bra .
De var utmärkta .
Han knackade på dörren och väntade .
Du borde gå till en läkare .
Liisa ryckte på axlarna .
Liisa försökte se snäll och menlös ut .
Markku suckade av lättnad .
Lägenheten bestod bara av ett enda rum .
Jag känner igen dig .
Pojken befann sig i en kvistig situation .
Är du inte riktigt klok ?
Just då ringde telefonen .
Markku är en ganska vanlig typ .
Det blev tyst i rummet .
Gubben tog fram sin fickalmanacka och bläddrade i den .
På golvet stod två par skor .
Det tog Liisa och Markku en kvart att komma dit .
Alla mina ankor simmar på sjön .
Du har fått det du ville , lämna mig ifred nu .
Tom är inte lång .
Välkommen tillbaka .
Vi har saknat dig !
Hon försöker begå självmord .
Varför i helvete lever du såhär , Tom ?
Tvätta dina händer .
Vi säljer skor .
Mary är en väldigt söt tjej .
Jag är gravid .
Kvinnan är naken .
Mannen rev sig på hakan och funderade på vad han skulle göra .
Han är rädd för katter .
Jag behöver en bil .
Hon förklarade ett skämt .
Han varnade dig .
Hon varnade dig .
Du är en idiot !
Min bror slog igen dörren med en smäll efter sig när han gick .
Liisa ruskade på huvudet .
Min far visste inte vad han skulle säga .
Jag känner mig vissen .
Jag har frågor .
Du sa till honom .
Sätt i ett mynt .
Det är ovanligt .
Jag gillar inte klassisk musik .
Jag måste lära mig ett språk .
Jag kommer att följa dig .
Är du rädd för höjder ?
Behöver du något ?
Jag behöver en bok att läsa .
Jag dricker vatten i köket .
Han kan ruttna i helvetet .
När blir det klart ?
Han ger ut böcker i Italien .
Jag vill skriva en bok .
Min lycka beror på dig .
Köpte du läkemedlet ?
De kallar den här planeten " Jord " .
Jag gillar mörk choklad .
Jag gillar katter mer än hundar .
Jag vet vad som gör mig lycklig .
Jag vet ingenting om det .
Människan uppfann atombomben , men ingen mus hade någonsin kommit på idén att konstruera en musfälla !
Storebror ser dig .
Jag vill inte göra några misstag .
Jag gör det om de betalar mig .
Vad är det ? frågade Tony .
Emet gillar inte den kvinnan .
Hej allihopa !
Du kan skriva på vilket språk du vill .
På Tatoeba är alla språk jämlika .
Markku verkade glatt överraskad .
Jag behöver inte uppehålsstillåtelse , för att jag är från Island .
Vi vill att regeringen ska tjäna hela befolkningen .
Vi vill att regeringen ska tjäna hela nationen .
Emet ogillar den där kvinnan .
Behöver ni någonting ?
Sjärnorna ser mycket vackra ut i kväll .
Detta är ett misstag .
Jag vill vara fri .
Jag vill inte begå några misstag .
Du har fått det du ville .
Lämna mig i fred nu .
Varför i helvete lever du så här , Tom ?
Studera de här meningarna .
Hon kan vare sig läsa eller skriva .
Där blev han anfallen av rebellerna .
Hon kan varken läsa eller skriva .
Jag kan rekommendera ett bra hotell .
Hon kan inte vare sig läsa eller skriva .
Vilka är dina fritidsintressen ?
On jest gruby .
Ingen knackar på min dörr .
Hur ser en vanlig dag ut för dig ?
Jag läser inte så många böcker som jag gjorde tidigare .
Förstår du vad jag menar ?
Det lever många hästar runt omkring mig .
Hur många hästar finns det i Sverige ?
Vi hjälpte dem .
Vi såg inget konstigt .
Det är inte längre klart var samhället slutar och var det privat kommersiella börjar .
Betty gick till havet i går .
Jag tycker om en skymning .
Vi har ingen dotter .
Min syster leker med dockan .
Fanns inga moln på himlen .
Upp med händerna !
Detta är ett rån .
Jag gör mitt bästa .
Man kan inte leva utan vatten .
Blomman är röd .
Han lagade en middag för henne .
Det här är mitt rum .
Jag lovar att säga till om jag ser något passande .
Kaffe och cigaretter .
Himlen och helvetet existerar i mans hjärtor .
Jag talar lite franska .
Stäng fönstret .
Öppna fönstret !
Öppna fönstret .
Han lärde sig att skriva siffror innan han kom till skolan .
Jag går till kyrkan .
Hon kan spela gitarr .
Tom är en kommunist .
Jag kan inte hjälpa dig .
Åker du med tåget eller bilen ?
Jag läser boken , medan jag äter .
Du får inte läsa , medan du äter .
Jag brukade inte röka .
Det är en film som alla borde se .
Vad kostar det ?
Jag har klardrömmar .
Min bror är väldigt lång .
Jag ser att du verkligen är en kåtbock ...
Ner på knä och slick min våta fitta !
Hädanefter är du min lydiga sexleksak .
Min lilla syster ockuperade mitt rum .
Jag är skild .
Tror du att han är död ?
Är han död ?
Tom har en ko .
Jag kan inte hjälpa er .
Solenergitekniken är kostnadseffektiv nuförtiden .
Jag vet var han är .
Hon bytte ämnet .
Jag måste åka till Danmark i morgon .
Vad är vi skyldiga ?
Vi var tvungna att gå till fots .
Jag tar hand om det .
Telefonen är trasig .
Det beror på stolens storlek .
Ditt förslag är lite extremt .
Tänker du ligga i sängen hela dagen , eller ?
Hur lärde du känna henne ?
Matematik är som kärlek – ett enkelt koncept , men det kan bli komplicerat .
Det är där jag kommer att vara .
Pojkarna och flickorna leker i trädgården .
Min engelsklärare rekommenderade mig att läsa dessa böcker .
Min engelsklärare rekommenderade mig att läsa de här böckerna .
Skulle ni kunna ta en titt på mitt första inlägg och berätta vad ni tycker om det ?
Tom tog bussen till skolan .
Tom tog en penna och började skriva .
Tom tog ut en penna och började skriva .
Tom tog av sig rocken eftersom det var för varmt för att ha den på sig .
Tom tog av sig rocken och kastade den på golvet .
Tom tog av sig sin rock och sina handskar .
Tom tog av sig sina kläder och gick in i duschen .
Hon är mycket vacker .
Att förstå dig är verkligen riktigt svårt .
Jämfört med hans far är han väldigt ytlig .
" Varför vill du så gärna dö ? "
" Varför vill du så gärna leva ? "
Det är verkligen riktigt svårt att förstå dig .
Vid slutet av den här månaden kommer antalet arbetande människor i den här staden att överstiga 1000 .
Det här är den högsta byggnad jag någonsin sett .
Tom tog av sig kläderna och gick in i duschen .
Detta är den högsta byggnad som jag någonsin har sett .
Detta är den högsta byggnad jag någonsin sett .
Detta är den högsta byggnad som jag någonsin sett .
Detta är den högsta byggnad jag någonsin har sett .
Det här är den högsta byggnad som jag någonsin sett .
Det här är den högsta byggnad jag någonsin har sett .
Tom tog av sig rocken och handskarna .
Tom tog fram en penna och började skriva .
Jag hjälpte henne med att hänga upp bilden på väggen .
Var är dina barn ?
Vad är växelkursen ?
Jag är mycket trött .
Jag är i Ryssland .
Han är mycket lång .
Har du varit i Kyoto ?
Jag såg henne igår .
Dörren är öppen .
Jag såg henne i går .
Han är mycket lång .
Var är era barn ?
Gillar du insekter ?
